`timescale 1 ns / 1 ns
module bandpass_filter_tb;

	parameter PERIOD = 4;

	reg clk, clk_en, rst_n;

	reg  signed [17:0] filter_in;
	wire signed [17:0] filter_out;

	reg  signed [17:0] filter_in_data_log_force [0:3148];
	reg  signed [17:0] filter_out_expected [0:3148];
	
	integer error, i, j;

	bandpass_filter b_filt 	(.i_clk(clk),
							 .i_clk_en(clk_en),
							 .i_rst_n(rst_n),
							 .i_data(filter_in),
							 .o_data(filter_out)
							 );

	initial begin
		clk = 0;
		forever #(PERIOD/2) clk = ~clk;
	end // initial

	initial begin
		error = 0;
		rst_n = 0;
		@(negedge clk);
		rst_n = 1;
		clk_en = 1;
		@(negedge clk);
		for (i=0; i<3149; i=i+1) begin 
			filter_in = filter_in_data_log_force[i];
			repeat(16) @(negedge clk);
		end
		
	end
	initial begin
		for (j=0; j<3149; j=j+1) begin 
			if (j==0) begin 
				repeat(33) @(negedge clk);
				if(filter_out !== filter_out_expected[j]) begin
					error = error + 1;
					$display("Error at time %d. Filter_out_real:%d Filter_out_expected[%d]:%d",
						$time, filter_out, j, filter_out_expected[j]);
				end
			end
			else begin
				repeat(16) @(posedge clk);
				@(negedge clk);
				if(filter_out !== filter_out_expected[j]) begin
					error = error + 1;
					$display("Error at time %d. Filter_out_real:%d Filter_out_expected[%d]:%d",
						$time, filter_out, j, filter_out_expected[j]);
				end
			end
		end
		if(error == 0)	$display("Test completed succesfully");
		else $display("Failed. Number of errors: %d",error);
		$finish;
	end
	initial begin
			
	 filter_in_data_log_force[   0] <= 18'h1ffff;
	 filter_in_data_log_force[   1] <= 18'h00000;
	 filter_in_data_log_force[   2] <= 18'h00000;
	 filter_in_data_log_force[   3] <= 18'h00000;
	 filter_in_data_log_force[   4] <= 18'h00000;
	 filter_in_data_log_force[   5] <= 18'h00000;
	 filter_in_data_log_force[   6] <= 18'h00000;
	 filter_in_data_log_force[   7] <= 18'h00000;
	 filter_in_data_log_force[   8] <= 18'h00000;
	 filter_in_data_log_force[   9] <= 18'h00000;
	 filter_in_data_log_force[  10] <= 18'h00000;
	 filter_in_data_log_force[  11] <= 18'h00000;
	 filter_in_data_log_force[  12] <= 18'h00000;
	 filter_in_data_log_force[  13] <= 18'h00000;
	 filter_in_data_log_force[  14] <= 18'h00000;
	 filter_in_data_log_force[  15] <= 18'h00000;
	 filter_in_data_log_force[  16] <= 18'h00000;
	 filter_in_data_log_force[  17] <= 18'h00000;
	 filter_in_data_log_force[  18] <= 18'h00000;
	 filter_in_data_log_force[  19] <= 18'h00000;
	 filter_in_data_log_force[  20] <= 18'h00000;
	 filter_in_data_log_force[  21] <= 18'h00000;
	 filter_in_data_log_force[  22] <= 18'h00000;
	 filter_in_data_log_force[  23] <= 18'h1ffff;
	 filter_in_data_log_force[  24] <= 18'h1ffff;
	 filter_in_data_log_force[  25] <= 18'h1ffff;
	 filter_in_data_log_force[  26] <= 18'h1ffff;
	 filter_in_data_log_force[  27] <= 18'h1ffff;
	 filter_in_data_log_force[  28] <= 18'h1ffff;
	 filter_in_data_log_force[  29] <= 18'h1ffff;
	 filter_in_data_log_force[  30] <= 18'h1ffff;
	 filter_in_data_log_force[  31] <= 18'h1ffff;
	 filter_in_data_log_force[  32] <= 18'h1ffff;
	 filter_in_data_log_force[  33] <= 18'h00000;
	 filter_in_data_log_force[  34] <= 18'h00000;
	 filter_in_data_log_force[  35] <= 18'h00000;
	 filter_in_data_log_force[  36] <= 18'h00000;
	 filter_in_data_log_force[  37] <= 18'h00000;
	 filter_in_data_log_force[  38] <= 18'h00000;
	 filter_in_data_log_force[  39] <= 18'h00000;
	 filter_in_data_log_force[  40] <= 18'h00000;
	 filter_in_data_log_force[  41] <= 18'h00000;
	 filter_in_data_log_force[  42] <= 18'h00000;
	 filter_in_data_log_force[  43] <= 18'h00000;
	 filter_in_data_log_force[  44] <= 18'h20000;
	 filter_in_data_log_force[  45] <= 18'h20100;
	 filter_in_data_log_force[  46] <= 18'h20201;
	 filter_in_data_log_force[  47] <= 18'h20301;
	 filter_in_data_log_force[  48] <= 18'h20401;
	 filter_in_data_log_force[  49] <= 18'h20501;
	 filter_in_data_log_force[  50] <= 18'h20602;
	 filter_in_data_log_force[  51] <= 18'h20702;
	 filter_in_data_log_force[  52] <= 18'h20802;
	 filter_in_data_log_force[  53] <= 18'h20902;
	 filter_in_data_log_force[  54] <= 18'h20a03;
	 filter_in_data_log_force[  55] <= 18'h20b03;
	 filter_in_data_log_force[  56] <= 18'h20c03;
	 filter_in_data_log_force[  57] <= 18'h20d03;
	 filter_in_data_log_force[  58] <= 18'h20e04;
	 filter_in_data_log_force[  59] <= 18'h20f04;
	 filter_in_data_log_force[  60] <= 18'h21004;
	 filter_in_data_log_force[  61] <= 18'h21104;
	 filter_in_data_log_force[  62] <= 18'h21205;
	 filter_in_data_log_force[  63] <= 18'h21305;
	 filter_in_data_log_force[  64] <= 18'h21405;
	 filter_in_data_log_force[  65] <= 18'h21505;
	 filter_in_data_log_force[  66] <= 18'h21606;
	 filter_in_data_log_force[  67] <= 18'h21706;
	 filter_in_data_log_force[  68] <= 18'h21806;
	 filter_in_data_log_force[  69] <= 18'h21906;
	 filter_in_data_log_force[  70] <= 18'h21a07;
	 filter_in_data_log_force[  71] <= 18'h21b07;
	 filter_in_data_log_force[  72] <= 18'h21c07;
	 filter_in_data_log_force[  73] <= 18'h21d07;
	 filter_in_data_log_force[  74] <= 18'h21e08;
	 filter_in_data_log_force[  75] <= 18'h21f08;
	 filter_in_data_log_force[  76] <= 18'h22008;
	 filter_in_data_log_force[  77] <= 18'h22108;
	 filter_in_data_log_force[  78] <= 18'h22209;
	 filter_in_data_log_force[  79] <= 18'h22309;
	 filter_in_data_log_force[  80] <= 18'h22409;
	 filter_in_data_log_force[  81] <= 18'h22509;
	 filter_in_data_log_force[  82] <= 18'h2260a;
	 filter_in_data_log_force[  83] <= 18'h2270a;
	 filter_in_data_log_force[  84] <= 18'h2280a;
	 filter_in_data_log_force[  85] <= 18'h2290a;
	 filter_in_data_log_force[  86] <= 18'h22a0b;
	 filter_in_data_log_force[  87] <= 18'h22b0b;
	 filter_in_data_log_force[  88] <= 18'h22c0b;
	 filter_in_data_log_force[  89] <= 18'h22d0b;
	 filter_in_data_log_force[  90] <= 18'h22e0c;
	 filter_in_data_log_force[  91] <= 18'h22f0c;
	 filter_in_data_log_force[  92] <= 18'h2300c;
	 filter_in_data_log_force[  93] <= 18'h2310c;
	 filter_in_data_log_force[  94] <= 18'h2320d;
	 filter_in_data_log_force[  95] <= 18'h2330d;
	 filter_in_data_log_force[  96] <= 18'h2340d;
	 filter_in_data_log_force[  97] <= 18'h2350d;
	 filter_in_data_log_force[  98] <= 18'h2360e;
	 filter_in_data_log_force[  99] <= 18'h2370e;
	 filter_in_data_log_force[ 100] <= 18'h2380e;
	 filter_in_data_log_force[ 101] <= 18'h2390e;
	 filter_in_data_log_force[ 102] <= 18'h23a0f;
	 filter_in_data_log_force[ 103] <= 18'h23b0f;
	 filter_in_data_log_force[ 104] <= 18'h23c0f;
	 filter_in_data_log_force[ 105] <= 18'h23d0f;
	 filter_in_data_log_force[ 106] <= 18'h23e10;
	 filter_in_data_log_force[ 107] <= 18'h23f10;
	 filter_in_data_log_force[ 108] <= 18'h24010;
	 filter_in_data_log_force[ 109] <= 18'h24110;
	 filter_in_data_log_force[ 110] <= 18'h24211;
	 filter_in_data_log_force[ 111] <= 18'h24311;
	 filter_in_data_log_force[ 112] <= 18'h24411;
	 filter_in_data_log_force[ 113] <= 18'h24511;
	 filter_in_data_log_force[ 114] <= 18'h24612;
	 filter_in_data_log_force[ 115] <= 18'h24712;
	 filter_in_data_log_force[ 116] <= 18'h24812;
	 filter_in_data_log_force[ 117] <= 18'h24912;
	 filter_in_data_log_force[ 118] <= 18'h24a13;
	 filter_in_data_log_force[ 119] <= 18'h24b13;
	 filter_in_data_log_force[ 120] <= 18'h24c13;
	 filter_in_data_log_force[ 121] <= 18'h24d13;
	 filter_in_data_log_force[ 122] <= 18'h24e14;
	 filter_in_data_log_force[ 123] <= 18'h24f14;
	 filter_in_data_log_force[ 124] <= 18'h25014;
	 filter_in_data_log_force[ 125] <= 18'h25114;
	 filter_in_data_log_force[ 126] <= 18'h25215;
	 filter_in_data_log_force[ 127] <= 18'h25315;
	 filter_in_data_log_force[ 128] <= 18'h25415;
	 filter_in_data_log_force[ 129] <= 18'h25515;
	 filter_in_data_log_force[ 130] <= 18'h25616;
	 filter_in_data_log_force[ 131] <= 18'h25716;
	 filter_in_data_log_force[ 132] <= 18'h25816;
	 filter_in_data_log_force[ 133] <= 18'h25916;
	 filter_in_data_log_force[ 134] <= 18'h25a17;
	 filter_in_data_log_force[ 135] <= 18'h25b17;
	 filter_in_data_log_force[ 136] <= 18'h25c17;
	 filter_in_data_log_force[ 137] <= 18'h25d17;
	 filter_in_data_log_force[ 138] <= 18'h25e18;
	 filter_in_data_log_force[ 139] <= 18'h25f18;
	 filter_in_data_log_force[ 140] <= 18'h26018;
	 filter_in_data_log_force[ 141] <= 18'h26118;
	 filter_in_data_log_force[ 142] <= 18'h26219;
	 filter_in_data_log_force[ 143] <= 18'h26319;
	 filter_in_data_log_force[ 144] <= 18'h26419;
	 filter_in_data_log_force[ 145] <= 18'h26519;
	 filter_in_data_log_force[ 146] <= 18'h2661a;
	 filter_in_data_log_force[ 147] <= 18'h2671a;
	 filter_in_data_log_force[ 148] <= 18'h2681a;
	 filter_in_data_log_force[ 149] <= 18'h2691a;
	 filter_in_data_log_force[ 150] <= 18'h26a1b;
	 filter_in_data_log_force[ 151] <= 18'h26b1b;
	 filter_in_data_log_force[ 152] <= 18'h26c1b;
	 filter_in_data_log_force[ 153] <= 18'h26d1b;
	 filter_in_data_log_force[ 154] <= 18'h26e1c;
	 filter_in_data_log_force[ 155] <= 18'h26f1c;
	 filter_in_data_log_force[ 156] <= 18'h2701c;
	 filter_in_data_log_force[ 157] <= 18'h2711c;
	 filter_in_data_log_force[ 158] <= 18'h2721d;
	 filter_in_data_log_force[ 159] <= 18'h2731d;
	 filter_in_data_log_force[ 160] <= 18'h2741d;
	 filter_in_data_log_force[ 161] <= 18'h2751d;
	 filter_in_data_log_force[ 162] <= 18'h2761e;
	 filter_in_data_log_force[ 163] <= 18'h2771e;
	 filter_in_data_log_force[ 164] <= 18'h2781e;
	 filter_in_data_log_force[ 165] <= 18'h2791e;
	 filter_in_data_log_force[ 166] <= 18'h27a1f;
	 filter_in_data_log_force[ 167] <= 18'h27b1f;
	 filter_in_data_log_force[ 168] <= 18'h27c1f;
	 filter_in_data_log_force[ 169] <= 18'h27d1f;
	 filter_in_data_log_force[ 170] <= 18'h27e20;
	 filter_in_data_log_force[ 171] <= 18'h27f20;
	 filter_in_data_log_force[ 172] <= 18'h28020;
	 filter_in_data_log_force[ 173] <= 18'h28120;
	 filter_in_data_log_force[ 174] <= 18'h28221;
	 filter_in_data_log_force[ 175] <= 18'h28321;
	 filter_in_data_log_force[ 176] <= 18'h28421;
	 filter_in_data_log_force[ 177] <= 18'h28521;
	 filter_in_data_log_force[ 178] <= 18'h28622;
	 filter_in_data_log_force[ 179] <= 18'h28722;
	 filter_in_data_log_force[ 180] <= 18'h28822;
	 filter_in_data_log_force[ 181] <= 18'h28922;
	 filter_in_data_log_force[ 182] <= 18'h28a23;
	 filter_in_data_log_force[ 183] <= 18'h28b23;
	 filter_in_data_log_force[ 184] <= 18'h28c23;
	 filter_in_data_log_force[ 185] <= 18'h28d23;
	 filter_in_data_log_force[ 186] <= 18'h28e24;
	 filter_in_data_log_force[ 187] <= 18'h28f24;
	 filter_in_data_log_force[ 188] <= 18'h29024;
	 filter_in_data_log_force[ 189] <= 18'h29124;
	 filter_in_data_log_force[ 190] <= 18'h29225;
	 filter_in_data_log_force[ 191] <= 18'h29325;
	 filter_in_data_log_force[ 192] <= 18'h29425;
	 filter_in_data_log_force[ 193] <= 18'h29525;
	 filter_in_data_log_force[ 194] <= 18'h29626;
	 filter_in_data_log_force[ 195] <= 18'h29726;
	 filter_in_data_log_force[ 196] <= 18'h29826;
	 filter_in_data_log_force[ 197] <= 18'h29926;
	 filter_in_data_log_force[ 198] <= 18'h29a27;
	 filter_in_data_log_force[ 199] <= 18'h29b27;
	 filter_in_data_log_force[ 200] <= 18'h29c27;
	 filter_in_data_log_force[ 201] <= 18'h29d27;
	 filter_in_data_log_force[ 202] <= 18'h29e28;
	 filter_in_data_log_force[ 203] <= 18'h29f28;
	 filter_in_data_log_force[ 204] <= 18'h2a028;
	 filter_in_data_log_force[ 205] <= 18'h2a128;
	 filter_in_data_log_force[ 206] <= 18'h2a229;
	 filter_in_data_log_force[ 207] <= 18'h2a329;
	 filter_in_data_log_force[ 208] <= 18'h2a429;
	 filter_in_data_log_force[ 209] <= 18'h2a529;
	 filter_in_data_log_force[ 210] <= 18'h2a62a;
	 filter_in_data_log_force[ 211] <= 18'h2a72a;
	 filter_in_data_log_force[ 212] <= 18'h2a82a;
	 filter_in_data_log_force[ 213] <= 18'h2a92a;
	 filter_in_data_log_force[ 214] <= 18'h2aa2b;
	 filter_in_data_log_force[ 215] <= 18'h2ab2b;
	 filter_in_data_log_force[ 216] <= 18'h2ac2b;
	 filter_in_data_log_force[ 217] <= 18'h2ad2b;
	 filter_in_data_log_force[ 218] <= 18'h2ae2c;
	 filter_in_data_log_force[ 219] <= 18'h2af2c;
	 filter_in_data_log_force[ 220] <= 18'h2b02c;
	 filter_in_data_log_force[ 221] <= 18'h2b12c;
	 filter_in_data_log_force[ 222] <= 18'h2b22d;
	 filter_in_data_log_force[ 223] <= 18'h2b32d;
	 filter_in_data_log_force[ 224] <= 18'h2b42d;
	 filter_in_data_log_force[ 225] <= 18'h2b52d;
	 filter_in_data_log_force[ 226] <= 18'h2b62e;
	 filter_in_data_log_force[ 227] <= 18'h2b72e;
	 filter_in_data_log_force[ 228] <= 18'h2b82e;
	 filter_in_data_log_force[ 229] <= 18'h2b92e;
	 filter_in_data_log_force[ 230] <= 18'h2ba2f;
	 filter_in_data_log_force[ 231] <= 18'h2bb2f;
	 filter_in_data_log_force[ 232] <= 18'h2bc2f;
	 filter_in_data_log_force[ 233] <= 18'h2bd2f;
	 filter_in_data_log_force[ 234] <= 18'h2be30;
	 filter_in_data_log_force[ 235] <= 18'h2bf30;
	 filter_in_data_log_force[ 236] <= 18'h2c030;
	 filter_in_data_log_force[ 237] <= 18'h2c130;
	 filter_in_data_log_force[ 238] <= 18'h2c231;
	 filter_in_data_log_force[ 239] <= 18'h2c331;
	 filter_in_data_log_force[ 240] <= 18'h2c431;
	 filter_in_data_log_force[ 241] <= 18'h2c531;
	 filter_in_data_log_force[ 242] <= 18'h2c632;
	 filter_in_data_log_force[ 243] <= 18'h2c732;
	 filter_in_data_log_force[ 244] <= 18'h2c832;
	 filter_in_data_log_force[ 245] <= 18'h2c932;
	 filter_in_data_log_force[ 246] <= 18'h2ca33;
	 filter_in_data_log_force[ 247] <= 18'h2cb33;
	 filter_in_data_log_force[ 248] <= 18'h2cc33;
	 filter_in_data_log_force[ 249] <= 18'h2cd33;
	 filter_in_data_log_force[ 250] <= 18'h2ce34;
	 filter_in_data_log_force[ 251] <= 18'h2cf34;
	 filter_in_data_log_force[ 252] <= 18'h2d034;
	 filter_in_data_log_force[ 253] <= 18'h2d134;
	 filter_in_data_log_force[ 254] <= 18'h2d235;
	 filter_in_data_log_force[ 255] <= 18'h2d335;
	 filter_in_data_log_force[ 256] <= 18'h2d435;
	 filter_in_data_log_force[ 257] <= 18'h2d535;
	 filter_in_data_log_force[ 258] <= 18'h2d636;
	 filter_in_data_log_force[ 259] <= 18'h2d736;
	 filter_in_data_log_force[ 260] <= 18'h2d836;
	 filter_in_data_log_force[ 261] <= 18'h2d936;
	 filter_in_data_log_force[ 262] <= 18'h2da37;
	 filter_in_data_log_force[ 263] <= 18'h2db37;
	 filter_in_data_log_force[ 264] <= 18'h2dc37;
	 filter_in_data_log_force[ 265] <= 18'h2dd37;
	 filter_in_data_log_force[ 266] <= 18'h2de38;
	 filter_in_data_log_force[ 267] <= 18'h2df38;
	 filter_in_data_log_force[ 268] <= 18'h2e038;
	 filter_in_data_log_force[ 269] <= 18'h2e138;
	 filter_in_data_log_force[ 270] <= 18'h2e239;
	 filter_in_data_log_force[ 271] <= 18'h2e339;
	 filter_in_data_log_force[ 272] <= 18'h2e439;
	 filter_in_data_log_force[ 273] <= 18'h2e539;
	 filter_in_data_log_force[ 274] <= 18'h2e63a;
	 filter_in_data_log_force[ 275] <= 18'h2e73a;
	 filter_in_data_log_force[ 276] <= 18'h2e83a;
	 filter_in_data_log_force[ 277] <= 18'h2e93a;
	 filter_in_data_log_force[ 278] <= 18'h2ea3b;
	 filter_in_data_log_force[ 279] <= 18'h2eb3b;
	 filter_in_data_log_force[ 280] <= 18'h2ec3b;
	 filter_in_data_log_force[ 281] <= 18'h2ed3b;
	 filter_in_data_log_force[ 282] <= 18'h2ee3c;
	 filter_in_data_log_force[ 283] <= 18'h2ef3c;
	 filter_in_data_log_force[ 284] <= 18'h2f03c;
	 filter_in_data_log_force[ 285] <= 18'h2f13c;
	 filter_in_data_log_force[ 286] <= 18'h2f23d;
	 filter_in_data_log_force[ 287] <= 18'h2f33d;
	 filter_in_data_log_force[ 288] <= 18'h2f43d;
	 filter_in_data_log_force[ 289] <= 18'h2f53d;
	 filter_in_data_log_force[ 290] <= 18'h2f63e;
	 filter_in_data_log_force[ 291] <= 18'h2f73e;
	 filter_in_data_log_force[ 292] <= 18'h2f83e;
	 filter_in_data_log_force[ 293] <= 18'h2f93e;
	 filter_in_data_log_force[ 294] <= 18'h2fa3f;
	 filter_in_data_log_force[ 295] <= 18'h2fb3f;
	 filter_in_data_log_force[ 296] <= 18'h2fc3f;
	 filter_in_data_log_force[ 297] <= 18'h2fd3f;
	 filter_in_data_log_force[ 298] <= 18'h2fe40;
	 filter_in_data_log_force[ 299] <= 18'h2ff40;
	 filter_in_data_log_force[ 300] <= 18'h30040;
	 filter_in_data_log_force[ 301] <= 18'h30140;
	 filter_in_data_log_force[ 302] <= 18'h30241;
	 filter_in_data_log_force[ 303] <= 18'h30341;
	 filter_in_data_log_force[ 304] <= 18'h30441;
	 filter_in_data_log_force[ 305] <= 18'h30541;
	 filter_in_data_log_force[ 306] <= 18'h30642;
	 filter_in_data_log_force[ 307] <= 18'h30742;
	 filter_in_data_log_force[ 308] <= 18'h30842;
	 filter_in_data_log_force[ 309] <= 18'h30942;
	 filter_in_data_log_force[ 310] <= 18'h30a43;
	 filter_in_data_log_force[ 311] <= 18'h30b43;
	 filter_in_data_log_force[ 312] <= 18'h30c43;
	 filter_in_data_log_force[ 313] <= 18'h30d43;
	 filter_in_data_log_force[ 314] <= 18'h30e44;
	 filter_in_data_log_force[ 315] <= 18'h30f44;
	 filter_in_data_log_force[ 316] <= 18'h31044;
	 filter_in_data_log_force[ 317] <= 18'h31144;
	 filter_in_data_log_force[ 318] <= 18'h31245;
	 filter_in_data_log_force[ 319] <= 18'h31345;
	 filter_in_data_log_force[ 320] <= 18'h31445;
	 filter_in_data_log_force[ 321] <= 18'h31545;
	 filter_in_data_log_force[ 322] <= 18'h31646;
	 filter_in_data_log_force[ 323] <= 18'h31746;
	 filter_in_data_log_force[ 324] <= 18'h31846;
	 filter_in_data_log_force[ 325] <= 18'h31946;
	 filter_in_data_log_force[ 326] <= 18'h31a47;
	 filter_in_data_log_force[ 327] <= 18'h31b47;
	 filter_in_data_log_force[ 328] <= 18'h31c47;
	 filter_in_data_log_force[ 329] <= 18'h31d47;
	 filter_in_data_log_force[ 330] <= 18'h31e48;
	 filter_in_data_log_force[ 331] <= 18'h31f48;
	 filter_in_data_log_force[ 332] <= 18'h32048;
	 filter_in_data_log_force[ 333] <= 18'h32148;
	 filter_in_data_log_force[ 334] <= 18'h32249;
	 filter_in_data_log_force[ 335] <= 18'h32349;
	 filter_in_data_log_force[ 336] <= 18'h32449;
	 filter_in_data_log_force[ 337] <= 18'h32549;
	 filter_in_data_log_force[ 338] <= 18'h3264a;
	 filter_in_data_log_force[ 339] <= 18'h3274a;
	 filter_in_data_log_force[ 340] <= 18'h3284a;
	 filter_in_data_log_force[ 341] <= 18'h3294a;
	 filter_in_data_log_force[ 342] <= 18'h32a4b;
	 filter_in_data_log_force[ 343] <= 18'h32b4b;
	 filter_in_data_log_force[ 344] <= 18'h32c4b;
	 filter_in_data_log_force[ 345] <= 18'h32d4b;
	 filter_in_data_log_force[ 346] <= 18'h32e4c;
	 filter_in_data_log_force[ 347] <= 18'h32f4c;
	 filter_in_data_log_force[ 348] <= 18'h3304c;
	 filter_in_data_log_force[ 349] <= 18'h3314c;
	 filter_in_data_log_force[ 350] <= 18'h3324d;
	 filter_in_data_log_force[ 351] <= 18'h3334d;
	 filter_in_data_log_force[ 352] <= 18'h3344d;
	 filter_in_data_log_force[ 353] <= 18'h3354d;
	 filter_in_data_log_force[ 354] <= 18'h3364e;
	 filter_in_data_log_force[ 355] <= 18'h3374e;
	 filter_in_data_log_force[ 356] <= 18'h3384e;
	 filter_in_data_log_force[ 357] <= 18'h3394e;
	 filter_in_data_log_force[ 358] <= 18'h33a4f;
	 filter_in_data_log_force[ 359] <= 18'h33b4f;
	 filter_in_data_log_force[ 360] <= 18'h33c4f;
	 filter_in_data_log_force[ 361] <= 18'h33d4f;
	 filter_in_data_log_force[ 362] <= 18'h33e50;
	 filter_in_data_log_force[ 363] <= 18'h33f50;
	 filter_in_data_log_force[ 364] <= 18'h34050;
	 filter_in_data_log_force[ 365] <= 18'h34150;
	 filter_in_data_log_force[ 366] <= 18'h34251;
	 filter_in_data_log_force[ 367] <= 18'h34351;
	 filter_in_data_log_force[ 368] <= 18'h34451;
	 filter_in_data_log_force[ 369] <= 18'h34551;
	 filter_in_data_log_force[ 370] <= 18'h34652;
	 filter_in_data_log_force[ 371] <= 18'h34752;
	 filter_in_data_log_force[ 372] <= 18'h34852;
	 filter_in_data_log_force[ 373] <= 18'h34952;
	 filter_in_data_log_force[ 374] <= 18'h34a53;
	 filter_in_data_log_force[ 375] <= 18'h34b53;
	 filter_in_data_log_force[ 376] <= 18'h34c53;
	 filter_in_data_log_force[ 377] <= 18'h34d53;
	 filter_in_data_log_force[ 378] <= 18'h34e54;
	 filter_in_data_log_force[ 379] <= 18'h34f54;
	 filter_in_data_log_force[ 380] <= 18'h35054;
	 filter_in_data_log_force[ 381] <= 18'h35154;
	 filter_in_data_log_force[ 382] <= 18'h35255;
	 filter_in_data_log_force[ 383] <= 18'h35355;
	 filter_in_data_log_force[ 384] <= 18'h35455;
	 filter_in_data_log_force[ 385] <= 18'h35555;
	 filter_in_data_log_force[ 386] <= 18'h35656;
	 filter_in_data_log_force[ 387] <= 18'h35756;
	 filter_in_data_log_force[ 388] <= 18'h35856;
	 filter_in_data_log_force[ 389] <= 18'h35956;
	 filter_in_data_log_force[ 390] <= 18'h35a57;
	 filter_in_data_log_force[ 391] <= 18'h35b57;
	 filter_in_data_log_force[ 392] <= 18'h35c57;
	 filter_in_data_log_force[ 393] <= 18'h35d57;
	 filter_in_data_log_force[ 394] <= 18'h35e58;
	 filter_in_data_log_force[ 395] <= 18'h35f58;
	 filter_in_data_log_force[ 396] <= 18'h36058;
	 filter_in_data_log_force[ 397] <= 18'h36158;
	 filter_in_data_log_force[ 398] <= 18'h36259;
	 filter_in_data_log_force[ 399] <= 18'h36359;
	 filter_in_data_log_force[ 400] <= 18'h36459;
	 filter_in_data_log_force[ 401] <= 18'h36559;
	 filter_in_data_log_force[ 402] <= 18'h3665a;
	 filter_in_data_log_force[ 403] <= 18'h3675a;
	 filter_in_data_log_force[ 404] <= 18'h3685a;
	 filter_in_data_log_force[ 405] <= 18'h3695a;
	 filter_in_data_log_force[ 406] <= 18'h36a5b;
	 filter_in_data_log_force[ 407] <= 18'h36b5b;
	 filter_in_data_log_force[ 408] <= 18'h36c5b;
	 filter_in_data_log_force[ 409] <= 18'h36d5b;
	 filter_in_data_log_force[ 410] <= 18'h36e5c;
	 filter_in_data_log_force[ 411] <= 18'h36f5c;
	 filter_in_data_log_force[ 412] <= 18'h3705c;
	 filter_in_data_log_force[ 413] <= 18'h3715c;
	 filter_in_data_log_force[ 414] <= 18'h3725d;
	 filter_in_data_log_force[ 415] <= 18'h3735d;
	 filter_in_data_log_force[ 416] <= 18'h3745d;
	 filter_in_data_log_force[ 417] <= 18'h3755d;
	 filter_in_data_log_force[ 418] <= 18'h3765e;
	 filter_in_data_log_force[ 419] <= 18'h3775e;
	 filter_in_data_log_force[ 420] <= 18'h3785e;
	 filter_in_data_log_force[ 421] <= 18'h3795e;
	 filter_in_data_log_force[ 422] <= 18'h37a5f;
	 filter_in_data_log_force[ 423] <= 18'h37b5f;
	 filter_in_data_log_force[ 424] <= 18'h37c5f;
	 filter_in_data_log_force[ 425] <= 18'h37d5f;
	 filter_in_data_log_force[ 426] <= 18'h37e60;
	 filter_in_data_log_force[ 427] <= 18'h37f60;
	 filter_in_data_log_force[ 428] <= 18'h38060;
	 filter_in_data_log_force[ 429] <= 18'h38160;
	 filter_in_data_log_force[ 430] <= 18'h38261;
	 filter_in_data_log_force[ 431] <= 18'h38361;
	 filter_in_data_log_force[ 432] <= 18'h38461;
	 filter_in_data_log_force[ 433] <= 18'h38561;
	 filter_in_data_log_force[ 434] <= 18'h38662;
	 filter_in_data_log_force[ 435] <= 18'h38762;
	 filter_in_data_log_force[ 436] <= 18'h38862;
	 filter_in_data_log_force[ 437] <= 18'h38962;
	 filter_in_data_log_force[ 438] <= 18'h38a63;
	 filter_in_data_log_force[ 439] <= 18'h38b63;
	 filter_in_data_log_force[ 440] <= 18'h38c63;
	 filter_in_data_log_force[ 441] <= 18'h38d63;
	 filter_in_data_log_force[ 442] <= 18'h38e64;
	 filter_in_data_log_force[ 443] <= 18'h38f64;
	 filter_in_data_log_force[ 444] <= 18'h39064;
	 filter_in_data_log_force[ 445] <= 18'h39164;
	 filter_in_data_log_force[ 446] <= 18'h39265;
	 filter_in_data_log_force[ 447] <= 18'h39365;
	 filter_in_data_log_force[ 448] <= 18'h39465;
	 filter_in_data_log_force[ 449] <= 18'h39565;
	 filter_in_data_log_force[ 450] <= 18'h39666;
	 filter_in_data_log_force[ 451] <= 18'h39766;
	 filter_in_data_log_force[ 452] <= 18'h39866;
	 filter_in_data_log_force[ 453] <= 18'h39966;
	 filter_in_data_log_force[ 454] <= 18'h39a67;
	 filter_in_data_log_force[ 455] <= 18'h39b67;
	 filter_in_data_log_force[ 456] <= 18'h39c67;
	 filter_in_data_log_force[ 457] <= 18'h39d67;
	 filter_in_data_log_force[ 458] <= 18'h39e68;
	 filter_in_data_log_force[ 459] <= 18'h39f68;
	 filter_in_data_log_force[ 460] <= 18'h3a068;
	 filter_in_data_log_force[ 461] <= 18'h3a168;
	 filter_in_data_log_force[ 462] <= 18'h3a269;
	 filter_in_data_log_force[ 463] <= 18'h3a369;
	 filter_in_data_log_force[ 464] <= 18'h3a469;
	 filter_in_data_log_force[ 465] <= 18'h3a569;
	 filter_in_data_log_force[ 466] <= 18'h3a66a;
	 filter_in_data_log_force[ 467] <= 18'h3a76a;
	 filter_in_data_log_force[ 468] <= 18'h3a86a;
	 filter_in_data_log_force[ 469] <= 18'h3a96a;
	 filter_in_data_log_force[ 470] <= 18'h3aa6b;
	 filter_in_data_log_force[ 471] <= 18'h3ab6b;
	 filter_in_data_log_force[ 472] <= 18'h3ac6b;
	 filter_in_data_log_force[ 473] <= 18'h3ad6b;
	 filter_in_data_log_force[ 474] <= 18'h3ae6c;
	 filter_in_data_log_force[ 475] <= 18'h3af6c;
	 filter_in_data_log_force[ 476] <= 18'h3b06c;
	 filter_in_data_log_force[ 477] <= 18'h3b16c;
	 filter_in_data_log_force[ 478] <= 18'h3b26d;
	 filter_in_data_log_force[ 479] <= 18'h3b36d;
	 filter_in_data_log_force[ 480] <= 18'h3b46d;
	 filter_in_data_log_force[ 481] <= 18'h3b56d;
	 filter_in_data_log_force[ 482] <= 18'h3b66e;
	 filter_in_data_log_force[ 483] <= 18'h3b76e;
	 filter_in_data_log_force[ 484] <= 18'h3b86e;
	 filter_in_data_log_force[ 485] <= 18'h3b96e;
	 filter_in_data_log_force[ 486] <= 18'h3ba6f;
	 filter_in_data_log_force[ 487] <= 18'h3bb6f;
	 filter_in_data_log_force[ 488] <= 18'h3bc6f;
	 filter_in_data_log_force[ 489] <= 18'h3bd6f;
	 filter_in_data_log_force[ 490] <= 18'h3be70;
	 filter_in_data_log_force[ 491] <= 18'h3bf70;
	 filter_in_data_log_force[ 492] <= 18'h3c070;
	 filter_in_data_log_force[ 493] <= 18'h3c170;
	 filter_in_data_log_force[ 494] <= 18'h3c271;
	 filter_in_data_log_force[ 495] <= 18'h3c371;
	 filter_in_data_log_force[ 496] <= 18'h3c471;
	 filter_in_data_log_force[ 497] <= 18'h3c571;
	 filter_in_data_log_force[ 498] <= 18'h3c672;
	 filter_in_data_log_force[ 499] <= 18'h3c772;
	 filter_in_data_log_force[ 500] <= 18'h3c872;
	 filter_in_data_log_force[ 501] <= 18'h3c972;
	 filter_in_data_log_force[ 502] <= 18'h3ca73;
	 filter_in_data_log_force[ 503] <= 18'h3cb73;
	 filter_in_data_log_force[ 504] <= 18'h3cc73;
	 filter_in_data_log_force[ 505] <= 18'h3cd73;
	 filter_in_data_log_force[ 506] <= 18'h3ce74;
	 filter_in_data_log_force[ 507] <= 18'h3cf74;
	 filter_in_data_log_force[ 508] <= 18'h3d074;
	 filter_in_data_log_force[ 509] <= 18'h3d174;
	 filter_in_data_log_force[ 510] <= 18'h3d275;
	 filter_in_data_log_force[ 511] <= 18'h3d375;
	 filter_in_data_log_force[ 512] <= 18'h3d475;
	 filter_in_data_log_force[ 513] <= 18'h3d575;
	 filter_in_data_log_force[ 514] <= 18'h3d676;
	 filter_in_data_log_force[ 515] <= 18'h3d776;
	 filter_in_data_log_force[ 516] <= 18'h3d876;
	 filter_in_data_log_force[ 517] <= 18'h3d976;
	 filter_in_data_log_force[ 518] <= 18'h3da77;
	 filter_in_data_log_force[ 519] <= 18'h3db77;
	 filter_in_data_log_force[ 520] <= 18'h3dc77;
	 filter_in_data_log_force[ 521] <= 18'h3dd77;
	 filter_in_data_log_force[ 522] <= 18'h3de78;
	 filter_in_data_log_force[ 523] <= 18'h3df78;
	 filter_in_data_log_force[ 524] <= 18'h3e078;
	 filter_in_data_log_force[ 525] <= 18'h3e178;
	 filter_in_data_log_force[ 526] <= 18'h3e279;
	 filter_in_data_log_force[ 527] <= 18'h3e379;
	 filter_in_data_log_force[ 528] <= 18'h3e479;
	 filter_in_data_log_force[ 529] <= 18'h3e579;
	 filter_in_data_log_force[ 530] <= 18'h3e67a;
	 filter_in_data_log_force[ 531] <= 18'h3e77a;
	 filter_in_data_log_force[ 532] <= 18'h3e87a;
	 filter_in_data_log_force[ 533] <= 18'h3e97a;
	 filter_in_data_log_force[ 534] <= 18'h3ea7b;
	 filter_in_data_log_force[ 535] <= 18'h3eb7b;
	 filter_in_data_log_force[ 536] <= 18'h3ec7b;
	 filter_in_data_log_force[ 537] <= 18'h3ed7b;
	 filter_in_data_log_force[ 538] <= 18'h3ee7c;
	 filter_in_data_log_force[ 539] <= 18'h3ef7c;
	 filter_in_data_log_force[ 540] <= 18'h3f07c;
	 filter_in_data_log_force[ 541] <= 18'h3f17c;
	 filter_in_data_log_force[ 542] <= 18'h3f27d;
	 filter_in_data_log_force[ 543] <= 18'h3f37d;
	 filter_in_data_log_force[ 544] <= 18'h3f47d;
	 filter_in_data_log_force[ 545] <= 18'h3f57d;
	 filter_in_data_log_force[ 546] <= 18'h3f67e;
	 filter_in_data_log_force[ 547] <= 18'h3f77e;
	 filter_in_data_log_force[ 548] <= 18'h3f87e;
	 filter_in_data_log_force[ 549] <= 18'h3f97e;
	 filter_in_data_log_force[ 550] <= 18'h3fa7f;
	 filter_in_data_log_force[ 551] <= 18'h3fb7f;
	 filter_in_data_log_force[ 552] <= 18'h3fc7f;
	 filter_in_data_log_force[ 553] <= 18'h3fd7f;
	 filter_in_data_log_force[ 554] <= 18'h3fe80;
	 filter_in_data_log_force[ 555] <= 18'h3ff80;
	 filter_in_data_log_force[ 556] <= 18'h00080;
	 filter_in_data_log_force[ 557] <= 18'h00180;
	 filter_in_data_log_force[ 558] <= 18'h00281;
	 filter_in_data_log_force[ 559] <= 18'h00381;
	 filter_in_data_log_force[ 560] <= 18'h00481;
	 filter_in_data_log_force[ 561] <= 18'h00581;
	 filter_in_data_log_force[ 562] <= 18'h00682;
	 filter_in_data_log_force[ 563] <= 18'h00782;
	 filter_in_data_log_force[ 564] <= 18'h00882;
	 filter_in_data_log_force[ 565] <= 18'h00982;
	 filter_in_data_log_force[ 566] <= 18'h00a83;
	 filter_in_data_log_force[ 567] <= 18'h00b83;
	 filter_in_data_log_force[ 568] <= 18'h00c83;
	 filter_in_data_log_force[ 569] <= 18'h00d83;
	 filter_in_data_log_force[ 570] <= 18'h00e84;
	 filter_in_data_log_force[ 571] <= 18'h00f84;
	 filter_in_data_log_force[ 572] <= 18'h01084;
	 filter_in_data_log_force[ 573] <= 18'h01184;
	 filter_in_data_log_force[ 574] <= 18'h01285;
	 filter_in_data_log_force[ 575] <= 18'h01385;
	 filter_in_data_log_force[ 576] <= 18'h01485;
	 filter_in_data_log_force[ 577] <= 18'h01585;
	 filter_in_data_log_force[ 578] <= 18'h01686;
	 filter_in_data_log_force[ 579] <= 18'h01786;
	 filter_in_data_log_force[ 580] <= 18'h01886;
	 filter_in_data_log_force[ 581] <= 18'h01986;
	 filter_in_data_log_force[ 582] <= 18'h01a87;
	 filter_in_data_log_force[ 583] <= 18'h01b87;
	 filter_in_data_log_force[ 584] <= 18'h01c87;
	 filter_in_data_log_force[ 585] <= 18'h01d87;
	 filter_in_data_log_force[ 586] <= 18'h01e88;
	 filter_in_data_log_force[ 587] <= 18'h01f88;
	 filter_in_data_log_force[ 588] <= 18'h02088;
	 filter_in_data_log_force[ 589] <= 18'h02188;
	 filter_in_data_log_force[ 590] <= 18'h02289;
	 filter_in_data_log_force[ 591] <= 18'h02389;
	 filter_in_data_log_force[ 592] <= 18'h02489;
	 filter_in_data_log_force[ 593] <= 18'h02589;
	 filter_in_data_log_force[ 594] <= 18'h0268a;
	 filter_in_data_log_force[ 595] <= 18'h0278a;
	 filter_in_data_log_force[ 596] <= 18'h0288a;
	 filter_in_data_log_force[ 597] <= 18'h0298a;
	 filter_in_data_log_force[ 598] <= 18'h02a8b;
	 filter_in_data_log_force[ 599] <= 18'h02b8b;
	 filter_in_data_log_force[ 600] <= 18'h02c8b;
	 filter_in_data_log_force[ 601] <= 18'h02d8b;
	 filter_in_data_log_force[ 602] <= 18'h02e8c;
	 filter_in_data_log_force[ 603] <= 18'h02f8c;
	 filter_in_data_log_force[ 604] <= 18'h0308c;
	 filter_in_data_log_force[ 605] <= 18'h0318c;
	 filter_in_data_log_force[ 606] <= 18'h0328d;
	 filter_in_data_log_force[ 607] <= 18'h0338d;
	 filter_in_data_log_force[ 608] <= 18'h0348d;
	 filter_in_data_log_force[ 609] <= 18'h0358d;
	 filter_in_data_log_force[ 610] <= 18'h0368e;
	 filter_in_data_log_force[ 611] <= 18'h0378e;
	 filter_in_data_log_force[ 612] <= 18'h0388e;
	 filter_in_data_log_force[ 613] <= 18'h0398e;
	 filter_in_data_log_force[ 614] <= 18'h03a8f;
	 filter_in_data_log_force[ 615] <= 18'h03b8f;
	 filter_in_data_log_force[ 616] <= 18'h03c8f;
	 filter_in_data_log_force[ 617] <= 18'h03d8f;
	 filter_in_data_log_force[ 618] <= 18'h03e90;
	 filter_in_data_log_force[ 619] <= 18'h03f90;
	 filter_in_data_log_force[ 620] <= 18'h04090;
	 filter_in_data_log_force[ 621] <= 18'h04190;
	 filter_in_data_log_force[ 622] <= 18'h04291;
	 filter_in_data_log_force[ 623] <= 18'h04391;
	 filter_in_data_log_force[ 624] <= 18'h04491;
	 filter_in_data_log_force[ 625] <= 18'h04591;
	 filter_in_data_log_force[ 626] <= 18'h04692;
	 filter_in_data_log_force[ 627] <= 18'h04792;
	 filter_in_data_log_force[ 628] <= 18'h04892;
	 filter_in_data_log_force[ 629] <= 18'h04992;
	 filter_in_data_log_force[ 630] <= 18'h04a93;
	 filter_in_data_log_force[ 631] <= 18'h04b93;
	 filter_in_data_log_force[ 632] <= 18'h04c93;
	 filter_in_data_log_force[ 633] <= 18'h04d93;
	 filter_in_data_log_force[ 634] <= 18'h04e94;
	 filter_in_data_log_force[ 635] <= 18'h04f94;
	 filter_in_data_log_force[ 636] <= 18'h05094;
	 filter_in_data_log_force[ 637] <= 18'h05194;
	 filter_in_data_log_force[ 638] <= 18'h05295;
	 filter_in_data_log_force[ 639] <= 18'h05395;
	 filter_in_data_log_force[ 640] <= 18'h05495;
	 filter_in_data_log_force[ 641] <= 18'h05595;
	 filter_in_data_log_force[ 642] <= 18'h05696;
	 filter_in_data_log_force[ 643] <= 18'h05796;
	 filter_in_data_log_force[ 644] <= 18'h05896;
	 filter_in_data_log_force[ 645] <= 18'h05996;
	 filter_in_data_log_force[ 646] <= 18'h05a97;
	 filter_in_data_log_force[ 647] <= 18'h05b97;
	 filter_in_data_log_force[ 648] <= 18'h05c97;
	 filter_in_data_log_force[ 649] <= 18'h05d97;
	 filter_in_data_log_force[ 650] <= 18'h05e98;
	 filter_in_data_log_force[ 651] <= 18'h05f98;
	 filter_in_data_log_force[ 652] <= 18'h06098;
	 filter_in_data_log_force[ 653] <= 18'h06198;
	 filter_in_data_log_force[ 654] <= 18'h06299;
	 filter_in_data_log_force[ 655] <= 18'h06399;
	 filter_in_data_log_force[ 656] <= 18'h06499;
	 filter_in_data_log_force[ 657] <= 18'h06599;
	 filter_in_data_log_force[ 658] <= 18'h0669a;
	 filter_in_data_log_force[ 659] <= 18'h0679a;
	 filter_in_data_log_force[ 660] <= 18'h0689a;
	 filter_in_data_log_force[ 661] <= 18'h0699a;
	 filter_in_data_log_force[ 662] <= 18'h06a9b;
	 filter_in_data_log_force[ 663] <= 18'h06b9b;
	 filter_in_data_log_force[ 664] <= 18'h06c9b;
	 filter_in_data_log_force[ 665] <= 18'h06d9b;
	 filter_in_data_log_force[ 666] <= 18'h06e9c;
	 filter_in_data_log_force[ 667] <= 18'h06f9c;
	 filter_in_data_log_force[ 668] <= 18'h0709c;
	 filter_in_data_log_force[ 669] <= 18'h0719c;
	 filter_in_data_log_force[ 670] <= 18'h0729d;
	 filter_in_data_log_force[ 671] <= 18'h0739d;
	 filter_in_data_log_force[ 672] <= 18'h0749d;
	 filter_in_data_log_force[ 673] <= 18'h0759d;
	 filter_in_data_log_force[ 674] <= 18'h0769e;
	 filter_in_data_log_force[ 675] <= 18'h0779e;
	 filter_in_data_log_force[ 676] <= 18'h0789e;
	 filter_in_data_log_force[ 677] <= 18'h0799e;
	 filter_in_data_log_force[ 678] <= 18'h07a9f;
	 filter_in_data_log_force[ 679] <= 18'h07b9f;
	 filter_in_data_log_force[ 680] <= 18'h07c9f;
	 filter_in_data_log_force[ 681] <= 18'h07d9f;
	 filter_in_data_log_force[ 682] <= 18'h07ea0;
	 filter_in_data_log_force[ 683] <= 18'h07fa0;
	 filter_in_data_log_force[ 684] <= 18'h080a0;
	 filter_in_data_log_force[ 685] <= 18'h081a0;
	 filter_in_data_log_force[ 686] <= 18'h082a1;
	 filter_in_data_log_force[ 687] <= 18'h083a1;
	 filter_in_data_log_force[ 688] <= 18'h084a1;
	 filter_in_data_log_force[ 689] <= 18'h085a1;
	 filter_in_data_log_force[ 690] <= 18'h086a2;
	 filter_in_data_log_force[ 691] <= 18'h087a2;
	 filter_in_data_log_force[ 692] <= 18'h088a2;
	 filter_in_data_log_force[ 693] <= 18'h089a2;
	 filter_in_data_log_force[ 694] <= 18'h08aa3;
	 filter_in_data_log_force[ 695] <= 18'h08ba3;
	 filter_in_data_log_force[ 696] <= 18'h08ca3;
	 filter_in_data_log_force[ 697] <= 18'h08da3;
	 filter_in_data_log_force[ 698] <= 18'h08ea4;
	 filter_in_data_log_force[ 699] <= 18'h08fa4;
	 filter_in_data_log_force[ 700] <= 18'h090a4;
	 filter_in_data_log_force[ 701] <= 18'h091a4;
	 filter_in_data_log_force[ 702] <= 18'h092a5;
	 filter_in_data_log_force[ 703] <= 18'h093a5;
	 filter_in_data_log_force[ 704] <= 18'h094a5;
	 filter_in_data_log_force[ 705] <= 18'h095a5;
	 filter_in_data_log_force[ 706] <= 18'h096a6;
	 filter_in_data_log_force[ 707] <= 18'h097a6;
	 filter_in_data_log_force[ 708] <= 18'h098a6;
	 filter_in_data_log_force[ 709] <= 18'h099a6;
	 filter_in_data_log_force[ 710] <= 18'h09aa7;
	 filter_in_data_log_force[ 711] <= 18'h09ba7;
	 filter_in_data_log_force[ 712] <= 18'h09ca7;
	 filter_in_data_log_force[ 713] <= 18'h09da7;
	 filter_in_data_log_force[ 714] <= 18'h09ea8;
	 filter_in_data_log_force[ 715] <= 18'h09fa8;
	 filter_in_data_log_force[ 716] <= 18'h0a0a8;
	 filter_in_data_log_force[ 717] <= 18'h0a1a8;
	 filter_in_data_log_force[ 718] <= 18'h0a2a9;
	 filter_in_data_log_force[ 719] <= 18'h0a3a9;
	 filter_in_data_log_force[ 720] <= 18'h0a4a9;
	 filter_in_data_log_force[ 721] <= 18'h0a5a9;
	 filter_in_data_log_force[ 722] <= 18'h0a6aa;
	 filter_in_data_log_force[ 723] <= 18'h0a7aa;
	 filter_in_data_log_force[ 724] <= 18'h0a8aa;
	 filter_in_data_log_force[ 725] <= 18'h0a9aa;
	 filter_in_data_log_force[ 726] <= 18'h0aaab;
	 filter_in_data_log_force[ 727] <= 18'h0abab;
	 filter_in_data_log_force[ 728] <= 18'h0acab;
	 filter_in_data_log_force[ 729] <= 18'h0adab;
	 filter_in_data_log_force[ 730] <= 18'h0aeac;
	 filter_in_data_log_force[ 731] <= 18'h0afac;
	 filter_in_data_log_force[ 732] <= 18'h0b0ac;
	 filter_in_data_log_force[ 733] <= 18'h0b1ac;
	 filter_in_data_log_force[ 734] <= 18'h0b2ad;
	 filter_in_data_log_force[ 735] <= 18'h0b3ad;
	 filter_in_data_log_force[ 736] <= 18'h0b4ad;
	 filter_in_data_log_force[ 737] <= 18'h0b5ad;
	 filter_in_data_log_force[ 738] <= 18'h0b6ae;
	 filter_in_data_log_force[ 739] <= 18'h0b7ae;
	 filter_in_data_log_force[ 740] <= 18'h0b8ae;
	 filter_in_data_log_force[ 741] <= 18'h0b9ae;
	 filter_in_data_log_force[ 742] <= 18'h0baaf;
	 filter_in_data_log_force[ 743] <= 18'h0bbaf;
	 filter_in_data_log_force[ 744] <= 18'h0bcaf;
	 filter_in_data_log_force[ 745] <= 18'h0bdaf;
	 filter_in_data_log_force[ 746] <= 18'h0beb0;
	 filter_in_data_log_force[ 747] <= 18'h0bfb0;
	 filter_in_data_log_force[ 748] <= 18'h0c0b0;
	 filter_in_data_log_force[ 749] <= 18'h0c1b0;
	 filter_in_data_log_force[ 750] <= 18'h0c2b1;
	 filter_in_data_log_force[ 751] <= 18'h0c3b1;
	 filter_in_data_log_force[ 752] <= 18'h0c4b1;
	 filter_in_data_log_force[ 753] <= 18'h0c5b1;
	 filter_in_data_log_force[ 754] <= 18'h0c6b2;
	 filter_in_data_log_force[ 755] <= 18'h0c7b2;
	 filter_in_data_log_force[ 756] <= 18'h0c8b2;
	 filter_in_data_log_force[ 757] <= 18'h0c9b2;
	 filter_in_data_log_force[ 758] <= 18'h0cab3;
	 filter_in_data_log_force[ 759] <= 18'h0cbb3;
	 filter_in_data_log_force[ 760] <= 18'h0ccb3;
	 filter_in_data_log_force[ 761] <= 18'h0cdb3;
	 filter_in_data_log_force[ 762] <= 18'h0ceb4;
	 filter_in_data_log_force[ 763] <= 18'h0cfb4;
	 filter_in_data_log_force[ 764] <= 18'h0d0b4;
	 filter_in_data_log_force[ 765] <= 18'h0d1b4;
	 filter_in_data_log_force[ 766] <= 18'h0d2b5;
	 filter_in_data_log_force[ 767] <= 18'h0d3b5;
	 filter_in_data_log_force[ 768] <= 18'h0d4b5;
	 filter_in_data_log_force[ 769] <= 18'h0d5b5;
	 filter_in_data_log_force[ 770] <= 18'h0d6b6;
	 filter_in_data_log_force[ 771] <= 18'h0d7b6;
	 filter_in_data_log_force[ 772] <= 18'h0d8b6;
	 filter_in_data_log_force[ 773] <= 18'h0d9b6;
	 filter_in_data_log_force[ 774] <= 18'h0dab7;
	 filter_in_data_log_force[ 775] <= 18'h0dbb7;
	 filter_in_data_log_force[ 776] <= 18'h0dcb7;
	 filter_in_data_log_force[ 777] <= 18'h0ddb7;
	 filter_in_data_log_force[ 778] <= 18'h0deb8;
	 filter_in_data_log_force[ 779] <= 18'h0dfb8;
	 filter_in_data_log_force[ 780] <= 18'h0e0b8;
	 filter_in_data_log_force[ 781] <= 18'h0e1b8;
	 filter_in_data_log_force[ 782] <= 18'h0e2b9;
	 filter_in_data_log_force[ 783] <= 18'h0e3b9;
	 filter_in_data_log_force[ 784] <= 18'h0e4b9;
	 filter_in_data_log_force[ 785] <= 18'h0e5b9;
	 filter_in_data_log_force[ 786] <= 18'h0e6ba;
	 filter_in_data_log_force[ 787] <= 18'h0e7ba;
	 filter_in_data_log_force[ 788] <= 18'h0e8ba;
	 filter_in_data_log_force[ 789] <= 18'h0e9ba;
	 filter_in_data_log_force[ 790] <= 18'h0eabb;
	 filter_in_data_log_force[ 791] <= 18'h0ebbb;
	 filter_in_data_log_force[ 792] <= 18'h0ecbb;
	 filter_in_data_log_force[ 793] <= 18'h0edbb;
	 filter_in_data_log_force[ 794] <= 18'h0eebc;
	 filter_in_data_log_force[ 795] <= 18'h0efbc;
	 filter_in_data_log_force[ 796] <= 18'h0f0bc;
	 filter_in_data_log_force[ 797] <= 18'h0f1bc;
	 filter_in_data_log_force[ 798] <= 18'h0f2bd;
	 filter_in_data_log_force[ 799] <= 18'h0f3bd;
	 filter_in_data_log_force[ 800] <= 18'h0f4bd;
	 filter_in_data_log_force[ 801] <= 18'h0f5bd;
	 filter_in_data_log_force[ 802] <= 18'h0f6be;
	 filter_in_data_log_force[ 803] <= 18'h0f7be;
	 filter_in_data_log_force[ 804] <= 18'h0f8be;
	 filter_in_data_log_force[ 805] <= 18'h0f9be;
	 filter_in_data_log_force[ 806] <= 18'h0fabf;
	 filter_in_data_log_force[ 807] <= 18'h0fbbf;
	 filter_in_data_log_force[ 808] <= 18'h0fcbf;
	 filter_in_data_log_force[ 809] <= 18'h0fdbf;
	 filter_in_data_log_force[ 810] <= 18'h0fec0;
	 filter_in_data_log_force[ 811] <= 18'h0ffc0;
	 filter_in_data_log_force[ 812] <= 18'h100c0;
	 filter_in_data_log_force[ 813] <= 18'h101c0;
	 filter_in_data_log_force[ 814] <= 18'h102c1;
	 filter_in_data_log_force[ 815] <= 18'h103c1;
	 filter_in_data_log_force[ 816] <= 18'h104c1;
	 filter_in_data_log_force[ 817] <= 18'h105c1;
	 filter_in_data_log_force[ 818] <= 18'h106c2;
	 filter_in_data_log_force[ 819] <= 18'h107c2;
	 filter_in_data_log_force[ 820] <= 18'h108c2;
	 filter_in_data_log_force[ 821] <= 18'h109c2;
	 filter_in_data_log_force[ 822] <= 18'h10ac3;
	 filter_in_data_log_force[ 823] <= 18'h10bc3;
	 filter_in_data_log_force[ 824] <= 18'h10cc3;
	 filter_in_data_log_force[ 825] <= 18'h10dc3;
	 filter_in_data_log_force[ 826] <= 18'h10ec4;
	 filter_in_data_log_force[ 827] <= 18'h10fc4;
	 filter_in_data_log_force[ 828] <= 18'h110c4;
	 filter_in_data_log_force[ 829] <= 18'h111c4;
	 filter_in_data_log_force[ 830] <= 18'h112c5;
	 filter_in_data_log_force[ 831] <= 18'h113c5;
	 filter_in_data_log_force[ 832] <= 18'h114c5;
	 filter_in_data_log_force[ 833] <= 18'h115c5;
	 filter_in_data_log_force[ 834] <= 18'h116c6;
	 filter_in_data_log_force[ 835] <= 18'h117c6;
	 filter_in_data_log_force[ 836] <= 18'h118c6;
	 filter_in_data_log_force[ 837] <= 18'h119c6;
	 filter_in_data_log_force[ 838] <= 18'h11ac7;
	 filter_in_data_log_force[ 839] <= 18'h11bc7;
	 filter_in_data_log_force[ 840] <= 18'h11cc7;
	 filter_in_data_log_force[ 841] <= 18'h11dc7;
	 filter_in_data_log_force[ 842] <= 18'h11ec8;
	 filter_in_data_log_force[ 843] <= 18'h11fc8;
	 filter_in_data_log_force[ 844] <= 18'h120c8;
	 filter_in_data_log_force[ 845] <= 18'h121c8;
	 filter_in_data_log_force[ 846] <= 18'h122c9;
	 filter_in_data_log_force[ 847] <= 18'h123c9;
	 filter_in_data_log_force[ 848] <= 18'h124c9;
	 filter_in_data_log_force[ 849] <= 18'h125c9;
	 filter_in_data_log_force[ 850] <= 18'h126ca;
	 filter_in_data_log_force[ 851] <= 18'h127ca;
	 filter_in_data_log_force[ 852] <= 18'h128ca;
	 filter_in_data_log_force[ 853] <= 18'h129ca;
	 filter_in_data_log_force[ 854] <= 18'h12acb;
	 filter_in_data_log_force[ 855] <= 18'h12bcb;
	 filter_in_data_log_force[ 856] <= 18'h12ccb;
	 filter_in_data_log_force[ 857] <= 18'h12dcb;
	 filter_in_data_log_force[ 858] <= 18'h12ecc;
	 filter_in_data_log_force[ 859] <= 18'h12fcc;
	 filter_in_data_log_force[ 860] <= 18'h130cc;
	 filter_in_data_log_force[ 861] <= 18'h131cc;
	 filter_in_data_log_force[ 862] <= 18'h132cd;
	 filter_in_data_log_force[ 863] <= 18'h133cd;
	 filter_in_data_log_force[ 864] <= 18'h134cd;
	 filter_in_data_log_force[ 865] <= 18'h135cd;
	 filter_in_data_log_force[ 866] <= 18'h136ce;
	 filter_in_data_log_force[ 867] <= 18'h137ce;
	 filter_in_data_log_force[ 868] <= 18'h138ce;
	 filter_in_data_log_force[ 869] <= 18'h139ce;
	 filter_in_data_log_force[ 870] <= 18'h13acf;
	 filter_in_data_log_force[ 871] <= 18'h13bcf;
	 filter_in_data_log_force[ 872] <= 18'h13ccf;
	 filter_in_data_log_force[ 873] <= 18'h13dcf;
	 filter_in_data_log_force[ 874] <= 18'h13ed0;
	 filter_in_data_log_force[ 875] <= 18'h13fd0;
	 filter_in_data_log_force[ 876] <= 18'h140d0;
	 filter_in_data_log_force[ 877] <= 18'h141d0;
	 filter_in_data_log_force[ 878] <= 18'h142d1;
	 filter_in_data_log_force[ 879] <= 18'h143d1;
	 filter_in_data_log_force[ 880] <= 18'h144d1;
	 filter_in_data_log_force[ 881] <= 18'h145d1;
	 filter_in_data_log_force[ 882] <= 18'h146d2;
	 filter_in_data_log_force[ 883] <= 18'h147d2;
	 filter_in_data_log_force[ 884] <= 18'h148d2;
	 filter_in_data_log_force[ 885] <= 18'h149d2;
	 filter_in_data_log_force[ 886] <= 18'h14ad3;
	 filter_in_data_log_force[ 887] <= 18'h14bd3;
	 filter_in_data_log_force[ 888] <= 18'h14cd3;
	 filter_in_data_log_force[ 889] <= 18'h14dd3;
	 filter_in_data_log_force[ 890] <= 18'h14ed4;
	 filter_in_data_log_force[ 891] <= 18'h14fd4;
	 filter_in_data_log_force[ 892] <= 18'h150d4;
	 filter_in_data_log_force[ 893] <= 18'h151d4;
	 filter_in_data_log_force[ 894] <= 18'h152d5;
	 filter_in_data_log_force[ 895] <= 18'h153d5;
	 filter_in_data_log_force[ 896] <= 18'h154d5;
	 filter_in_data_log_force[ 897] <= 18'h155d5;
	 filter_in_data_log_force[ 898] <= 18'h156d6;
	 filter_in_data_log_force[ 899] <= 18'h157d6;
	 filter_in_data_log_force[ 900] <= 18'h158d6;
	 filter_in_data_log_force[ 901] <= 18'h159d6;
	 filter_in_data_log_force[ 902] <= 18'h15ad7;
	 filter_in_data_log_force[ 903] <= 18'h15bd7;
	 filter_in_data_log_force[ 904] <= 18'h15cd7;
	 filter_in_data_log_force[ 905] <= 18'h15dd7;
	 filter_in_data_log_force[ 906] <= 18'h15ed8;
	 filter_in_data_log_force[ 907] <= 18'h15fd8;
	 filter_in_data_log_force[ 908] <= 18'h160d8;
	 filter_in_data_log_force[ 909] <= 18'h161d8;
	 filter_in_data_log_force[ 910] <= 18'h162d9;
	 filter_in_data_log_force[ 911] <= 18'h163d9;
	 filter_in_data_log_force[ 912] <= 18'h164d9;
	 filter_in_data_log_force[ 913] <= 18'h165d9;
	 filter_in_data_log_force[ 914] <= 18'h166da;
	 filter_in_data_log_force[ 915] <= 18'h167da;
	 filter_in_data_log_force[ 916] <= 18'h168da;
	 filter_in_data_log_force[ 917] <= 18'h169da;
	 filter_in_data_log_force[ 918] <= 18'h16adb;
	 filter_in_data_log_force[ 919] <= 18'h16bdb;
	 filter_in_data_log_force[ 920] <= 18'h16cdb;
	 filter_in_data_log_force[ 921] <= 18'h16ddb;
	 filter_in_data_log_force[ 922] <= 18'h16edc;
	 filter_in_data_log_force[ 923] <= 18'h16fdc;
	 filter_in_data_log_force[ 924] <= 18'h170dc;
	 filter_in_data_log_force[ 925] <= 18'h171dc;
	 filter_in_data_log_force[ 926] <= 18'h172dd;
	 filter_in_data_log_force[ 927] <= 18'h173dd;
	 filter_in_data_log_force[ 928] <= 18'h174dd;
	 filter_in_data_log_force[ 929] <= 18'h175dd;
	 filter_in_data_log_force[ 930] <= 18'h176de;
	 filter_in_data_log_force[ 931] <= 18'h177de;
	 filter_in_data_log_force[ 932] <= 18'h178de;
	 filter_in_data_log_force[ 933] <= 18'h179de;
	 filter_in_data_log_force[ 934] <= 18'h17adf;
	 filter_in_data_log_force[ 935] <= 18'h17bdf;
	 filter_in_data_log_force[ 936] <= 18'h17cdf;
	 filter_in_data_log_force[ 937] <= 18'h17ddf;
	 filter_in_data_log_force[ 938] <= 18'h17ee0;
	 filter_in_data_log_force[ 939] <= 18'h17fe0;
	 filter_in_data_log_force[ 940] <= 18'h180e0;
	 filter_in_data_log_force[ 941] <= 18'h181e0;
	 filter_in_data_log_force[ 942] <= 18'h182e1;
	 filter_in_data_log_force[ 943] <= 18'h183e1;
	 filter_in_data_log_force[ 944] <= 18'h184e1;
	 filter_in_data_log_force[ 945] <= 18'h185e1;
	 filter_in_data_log_force[ 946] <= 18'h186e2;
	 filter_in_data_log_force[ 947] <= 18'h187e2;
	 filter_in_data_log_force[ 948] <= 18'h188e2;
	 filter_in_data_log_force[ 949] <= 18'h189e2;
	 filter_in_data_log_force[ 950] <= 18'h18ae3;
	 filter_in_data_log_force[ 951] <= 18'h18be3;
	 filter_in_data_log_force[ 952] <= 18'h18ce3;
	 filter_in_data_log_force[ 953] <= 18'h18de3;
	 filter_in_data_log_force[ 954] <= 18'h18ee4;
	 filter_in_data_log_force[ 955] <= 18'h18fe4;
	 filter_in_data_log_force[ 956] <= 18'h190e4;
	 filter_in_data_log_force[ 957] <= 18'h191e4;
	 filter_in_data_log_force[ 958] <= 18'h192e5;
	 filter_in_data_log_force[ 959] <= 18'h193e5;
	 filter_in_data_log_force[ 960] <= 18'h194e5;
	 filter_in_data_log_force[ 961] <= 18'h195e5;
	 filter_in_data_log_force[ 962] <= 18'h196e6;
	 filter_in_data_log_force[ 963] <= 18'h197e6;
	 filter_in_data_log_force[ 964] <= 18'h198e6;
	 filter_in_data_log_force[ 965] <= 18'h199e6;
	 filter_in_data_log_force[ 966] <= 18'h19ae7;
	 filter_in_data_log_force[ 967] <= 18'h19be7;
	 filter_in_data_log_force[ 968] <= 18'h19ce7;
	 filter_in_data_log_force[ 969] <= 18'h19de7;
	 filter_in_data_log_force[ 970] <= 18'h19ee8;
	 filter_in_data_log_force[ 971] <= 18'h19fe8;
	 filter_in_data_log_force[ 972] <= 18'h1a0e8;
	 filter_in_data_log_force[ 973] <= 18'h1a1e8;
	 filter_in_data_log_force[ 974] <= 18'h1a2e9;
	 filter_in_data_log_force[ 975] <= 18'h1a3e9;
	 filter_in_data_log_force[ 976] <= 18'h1a4e9;
	 filter_in_data_log_force[ 977] <= 18'h1a5e9;
	 filter_in_data_log_force[ 978] <= 18'h1a6ea;
	 filter_in_data_log_force[ 979] <= 18'h1a7ea;
	 filter_in_data_log_force[ 980] <= 18'h1a8ea;
	 filter_in_data_log_force[ 981] <= 18'h1a9ea;
	 filter_in_data_log_force[ 982] <= 18'h1aaeb;
	 filter_in_data_log_force[ 983] <= 18'h1abeb;
	 filter_in_data_log_force[ 984] <= 18'h1aceb;
	 filter_in_data_log_force[ 985] <= 18'h1adeb;
	 filter_in_data_log_force[ 986] <= 18'h1aeec;
	 filter_in_data_log_force[ 987] <= 18'h1afec;
	 filter_in_data_log_force[ 988] <= 18'h1b0ec;
	 filter_in_data_log_force[ 989] <= 18'h1b1ec;
	 filter_in_data_log_force[ 990] <= 18'h1b2ed;
	 filter_in_data_log_force[ 991] <= 18'h1b3ed;
	 filter_in_data_log_force[ 992] <= 18'h1b4ed;
	 filter_in_data_log_force[ 993] <= 18'h1b5ed;
	 filter_in_data_log_force[ 994] <= 18'h1b6ee;
	 filter_in_data_log_force[ 995] <= 18'h1b7ee;
	 filter_in_data_log_force[ 996] <= 18'h1b8ee;
	 filter_in_data_log_force[ 997] <= 18'h1b9ee;
	 filter_in_data_log_force[ 998] <= 18'h1baef;
	 filter_in_data_log_force[ 999] <= 18'h1bbef;
	 filter_in_data_log_force[1000] <= 18'h1bcef;
	 filter_in_data_log_force[1001] <= 18'h1bdef;
	 filter_in_data_log_force[1002] <= 18'h1bef0;
	 filter_in_data_log_force[1003] <= 18'h1bff0;
	 filter_in_data_log_force[1004] <= 18'h1c0f0;
	 filter_in_data_log_force[1005] <= 18'h1c1f0;
	 filter_in_data_log_force[1006] <= 18'h1c2f1;
	 filter_in_data_log_force[1007] <= 18'h1c3f1;
	 filter_in_data_log_force[1008] <= 18'h1c4f1;
	 filter_in_data_log_force[1009] <= 18'h1c5f1;
	 filter_in_data_log_force[1010] <= 18'h1c6f2;
	 filter_in_data_log_force[1011] <= 18'h1c7f2;
	 filter_in_data_log_force[1012] <= 18'h1c8f2;
	 filter_in_data_log_force[1013] <= 18'h1c9f2;
	 filter_in_data_log_force[1014] <= 18'h1caf3;
	 filter_in_data_log_force[1015] <= 18'h1cbf3;
	 filter_in_data_log_force[1016] <= 18'h1ccf3;
	 filter_in_data_log_force[1017] <= 18'h1cdf3;
	 filter_in_data_log_force[1018] <= 18'h1cef4;
	 filter_in_data_log_force[1019] <= 18'h1cff4;
	 filter_in_data_log_force[1020] <= 18'h1d0f4;
	 filter_in_data_log_force[1021] <= 18'h1d1f4;
	 filter_in_data_log_force[1022] <= 18'h1d2f5;
	 filter_in_data_log_force[1023] <= 18'h1d3f5;
	 filter_in_data_log_force[1024] <= 18'h1d4f5;
	 filter_in_data_log_force[1025] <= 18'h1d5f5;
	 filter_in_data_log_force[1026] <= 18'h1d6f6;
	 filter_in_data_log_force[1027] <= 18'h1d7f6;
	 filter_in_data_log_force[1028] <= 18'h1d8f6;
	 filter_in_data_log_force[1029] <= 18'h1d9f6;
	 filter_in_data_log_force[1030] <= 18'h1daf7;
	 filter_in_data_log_force[1031] <= 18'h1dbf7;
	 filter_in_data_log_force[1032] <= 18'h1dcf7;
	 filter_in_data_log_force[1033] <= 18'h1ddf7;
	 filter_in_data_log_force[1034] <= 18'h1def8;
	 filter_in_data_log_force[1035] <= 18'h1dff8;
	 filter_in_data_log_force[1036] <= 18'h1e0f8;
	 filter_in_data_log_force[1037] <= 18'h1e1f8;
	 filter_in_data_log_force[1038] <= 18'h1e2f9;
	 filter_in_data_log_force[1039] <= 18'h1e3f9;
	 filter_in_data_log_force[1040] <= 18'h1e4f9;
	 filter_in_data_log_force[1041] <= 18'h1e5f9;
	 filter_in_data_log_force[1042] <= 18'h1e6fa;
	 filter_in_data_log_force[1043] <= 18'h1e7fa;
	 filter_in_data_log_force[1044] <= 18'h1e8fa;
	 filter_in_data_log_force[1045] <= 18'h1e9fa;
	 filter_in_data_log_force[1046] <= 18'h1eafb;
	 filter_in_data_log_force[1047] <= 18'h1ebfb;
	 filter_in_data_log_force[1048] <= 18'h1ecfb;
	 filter_in_data_log_force[1049] <= 18'h1edfb;
	 filter_in_data_log_force[1050] <= 18'h1eefc;
	 filter_in_data_log_force[1051] <= 18'h1effc;
	 filter_in_data_log_force[1052] <= 18'h1f0fc;
	 filter_in_data_log_force[1053] <= 18'h1f1fc;
	 filter_in_data_log_force[1054] <= 18'h1f2fd;
	 filter_in_data_log_force[1055] <= 18'h1f3fd;
	 filter_in_data_log_force[1056] <= 18'h1f4fd;
	 filter_in_data_log_force[1057] <= 18'h1f5fd;
	 filter_in_data_log_force[1058] <= 18'h1f6fe;
	 filter_in_data_log_force[1059] <= 18'h1f7fe;
	 filter_in_data_log_force[1060] <= 18'h1f8fe;
	 filter_in_data_log_force[1061] <= 18'h1f9fe;
	 filter_in_data_log_force[1062] <= 18'h1faff;
	 filter_in_data_log_force[1063] <= 18'h1fbff;
	 filter_in_data_log_force[1064] <= 18'h1fcff;
	 filter_in_data_log_force[1065] <= 18'h1fdff;
	 filter_in_data_log_force[1066] <= 18'h1ff00;
	 filter_in_data_log_force[1067] <= 18'h1ffff;
	 filter_in_data_log_force[1068] <= 18'h00000;
	 filter_in_data_log_force[1069] <= 18'h00000;
	 filter_in_data_log_force[1070] <= 18'h00000;
	 filter_in_data_log_force[1071] <= 18'h00000;
	 filter_in_data_log_force[1072] <= 18'h00000;
	 filter_in_data_log_force[1073] <= 18'h00000;
	 filter_in_data_log_force[1074] <= 18'h00000;
	 filter_in_data_log_force[1075] <= 18'h00000;
	 filter_in_data_log_force[1076] <= 18'h00000;
	 filter_in_data_log_force[1077] <= 18'h00000;
	 filter_in_data_log_force[1078] <= 18'h00000;
	 filter_in_data_log_force[1079] <= 18'h1ffff;
	 filter_in_data_log_force[1080] <= 18'h1ffff;
	 filter_in_data_log_force[1081] <= 18'h1fffe;
	 filter_in_data_log_force[1082] <= 18'h1fff4;
	 filter_in_data_log_force[1083] <= 18'h1ffda;
	 filter_in_data_log_force[1084] <= 18'h1ffa3;
	 filter_in_data_log_force[1085] <= 18'h1ff40;
	 filter_in_data_log_force[1086] <= 18'h1fe9c;
	 filter_in_data_log_force[1087] <= 18'h1fda1;
	 filter_in_data_log_force[1088] <= 18'h1fc34;
	 filter_in_data_log_force[1089] <= 18'h1fa37;
	 filter_in_data_log_force[1090] <= 18'h1f789;
	 filter_in_data_log_force[1091] <= 18'h1f407;
	 filter_in_data_log_force[1092] <= 18'h1ef88;
	 filter_in_data_log_force[1093] <= 18'h1e9e4;
	 filter_in_data_log_force[1094] <= 18'h1e2ef;
	 filter_in_data_log_force[1095] <= 18'h1da7a;
	 filter_in_data_log_force[1096] <= 18'h1d058;
	 filter_in_data_log_force[1097] <= 18'h1c458;
	 filter_in_data_log_force[1098] <= 18'h1b64c;
	 filter_in_data_log_force[1099] <= 18'h1a605;
	 filter_in_data_log_force[1100] <= 18'h19358;
	 filter_in_data_log_force[1101] <= 18'h17e1b;
	 filter_in_data_log_force[1102] <= 18'h1662c;
	 filter_in_data_log_force[1103] <= 18'h14b6c;
	 filter_in_data_log_force[1104] <= 18'h12dc6;
	 filter_in_data_log_force[1105] <= 18'h10d2c;
	 filter_in_data_log_force[1106] <= 18'h0e99f;
	 filter_in_data_log_force[1107] <= 18'h0c328;
	 filter_in_data_log_force[1108] <= 18'h099e4;
	 filter_in_data_log_force[1109] <= 18'h06dfc;
	 filter_in_data_log_force[1110] <= 18'h03fb0;
	 filter_in_data_log_force[1111] <= 18'h00f50;
	 filter_in_data_log_force[1112] <= 18'h3dd43;
	 filter_in_data_log_force[1113] <= 18'h3aa06;
	 filter_in_data_log_force[1114] <= 18'h3762d;
	 filter_in_data_log_force[1115] <= 18'h34261;
	 filter_in_data_log_force[1116] <= 18'h30f63;
	 filter_in_data_log_force[1117] <= 18'h2de05;
	 filter_in_data_log_force[1118] <= 18'h2af2e;
	 filter_in_data_log_force[1119] <= 18'h283d3;
	 filter_in_data_log_force[1120] <= 18'h25cf3;
	 filter_in_data_log_force[1121] <= 18'h23b91;
	 filter_in_data_log_force[1122] <= 18'h220b1;
	 filter_in_data_log_force[1123] <= 18'h20d4b;
	 filter_in_data_log_force[1124] <= 18'h20248;
	 filter_in_data_log_force[1125] <= 18'h20076;
	 filter_in_data_log_force[1126] <= 18'h2087f;
	 filter_in_data_log_force[1127] <= 18'h21ade;
	 filter_in_data_log_force[1128] <= 18'h237d5;
	 filter_in_data_log_force[1129] <= 18'h25f65;
	 filter_in_data_log_force[1130] <= 18'h29142;
	 filter_in_data_log_force[1131] <= 18'h2ccce;
	 filter_in_data_log_force[1132] <= 18'h31115;
	 filter_in_data_log_force[1133] <= 18'h35cc4;
	 filter_in_data_log_force[1134] <= 18'h3ae33;
	 filter_in_data_log_force[1135] <= 18'h0035d;
	 filter_in_data_log_force[1136] <= 18'h059f5;
	 filter_in_data_log_force[1137] <= 18'h0af66;
	 filter_in_data_log_force[1138] <= 18'h100f0;
	 filter_in_data_log_force[1139] <= 18'h14bb6;
	 filter_in_data_log_force[1140] <= 18'h18cd9;
	 filter_in_data_log_force[1141] <= 18'h1c19b;
	 filter_in_data_log_force[1142] <= 18'h1e77a;
	 filter_in_data_log_force[1143] <= 18'h1fc57;
	 filter_in_data_log_force[1144] <= 18'h1fe95;
	 filter_in_data_log_force[1145] <= 18'h1ed3b;
	 filter_in_data_log_force[1146] <= 18'h1c815;
	 filter_in_data_log_force[1147] <= 18'h18fc3;
	 filter_in_data_log_force[1148] <= 18'h145d1;
	 filter_in_data_log_force[1149] <= 18'h0ecb5;
	 filter_in_data_log_force[1150] <= 18'h087cb;
	 filter_in_data_log_force[1151] <= 18'h01b40;
	 filter_in_data_log_force[1152] <= 18'h3abef;
	 filter_in_data_log_force[1153] <= 18'h33f2c;
	 filter_in_data_log_force[1154] <= 18'h2da8b;
	 filter_in_data_log_force[1155] <= 18'h28393;
	 filter_in_data_log_force[1156] <= 18'h23f6a;
	 filter_in_data_log_force[1157] <= 18'h21284;
	 filter_in_data_log_force[1158] <= 18'h2004a;
	 filter_in_data_log_force[1159] <= 18'h20acd;
	 filter_in_data_log_force[1160] <= 18'h23288;
	 filter_in_data_log_force[1161] <= 18'h27633;
	 filter_in_data_log_force[1162] <= 18'h2d2af;
	 filter_in_data_log_force[1163] <= 18'h34315;
	 filter_in_data_log_force[1164] <= 18'h3c0e0;
	 filter_in_data_log_force[1165] <= 18'h04441;
	 filter_in_data_log_force[1166] <= 18'h0c491;
	 filter_in_data_log_force[1167] <= 18'h138da;
	 filter_in_data_log_force[1168] <= 18'h1987f;
	 filter_in_data_log_force[1169] <= 18'h1dbe8;
	 filter_in_data_log_force[1170] <= 18'h1fd29;
	 filter_in_data_log_force[1171] <= 18'h1f89e;
	 filter_in_data_log_force[1172] <= 18'h1cd63;
	 filter_in_data_log_force[1173] <= 18'h17d9a;
	 filter_in_data_log_force[1174] <= 18'h10e7f;
	 filter_in_data_log_force[1175] <= 18'h0882c;
	 filter_in_data_log_force[1176] <= 18'h3f523;
	 filter_in_data_log_force[1177] <= 18'h3618b;
	 filter_in_data_log_force[1178] <= 18'h2da3c;
	 filter_in_data_log_force[1179] <= 18'h26b9b;
	 filter_in_data_log_force[1180] <= 18'h2206d;
	 filter_in_data_log_force[1181] <= 18'h200b3;
	 filter_in_data_log_force[1182] <= 18'h210b5;
	 filter_in_data_log_force[1183] <= 18'h2504b;
	 filter_in_data_log_force[1184] <= 18'h2ba9f;
	 filter_in_data_log_force[1185] <= 18'h3464d;
	 filter_in_data_log_force[1186] <= 18'h3e615;
	 filter_in_data_log_force[1187] <= 18'h089fd;
	 filter_in_data_log_force[1188] <= 18'h120da;
	 filter_in_data_log_force[1189] <= 18'h19a1d;
	 filter_in_data_log_force[1190] <= 18'h1e7b5;
	 filter_in_data_log_force[1191] <= 18'h1ffd3;
	 filter_in_data_log_force[1192] <= 18'h1de4c;
	 filter_in_data_log_force[1193] <= 18'h18577;
	 filter_in_data_log_force[1194] <= 18'h0fe4c;
	 filter_in_data_log_force[1195] <= 18'h057b6;
	 filter_in_data_log_force[1196] <= 18'h3a51e;
	 filter_in_data_log_force[1197] <= 18'h2fc40;
	 filter_in_data_log_force[1198] <= 18'h2728f;
	 filter_in_data_log_force[1199] <= 18'h21a63;
	 filter_in_data_log_force[1200] <= 18'h2006a;
	 filter_in_data_log_force[1201] <= 18'h22998;
	 filter_in_data_log_force[1202] <= 18'h2920c;
	 filter_in_data_log_force[1203] <= 18'h32d15;
	 filter_in_data_log_force[1204] <= 18'h3e676;
	 filter_in_data_log_force[1205] <= 18'h0a4d7;
	 filter_in_data_log_force[1206] <= 18'h14d28;
	 filter_in_data_log_force[1207] <= 18'h1c67a;
	 filter_in_data_log_force[1208] <= 18'h1fdd7;
	 filter_in_data_log_force[1209] <= 18'h1e974;
	 filter_in_data_log_force[1210] <= 18'h18aac;
	 filter_in_data_log_force[1211] <= 18'h0ee6f;
	 filter_in_data_log_force[1212] <= 18'h02bcc;
	 filter_in_data_log_force[1213] <= 18'h360d4;
	 filter_in_data_log_force[1214] <= 18'h2ae0c;
	 filter_in_data_log_force[1215] <= 18'h2313a;
	 filter_in_data_log_force[1216] <= 18'h20040;
	 filter_in_data_log_force[1217] <= 18'h22501;
	 filter_in_data_log_force[1218] <= 18'h29b0b;
	 filter_in_data_log_force[1219] <= 18'h34fa8;
	 filter_in_data_log_force[1220] <= 18'h0246e;
	 filter_in_data_log_force[1221] <= 18'h0f425;
	 filter_in_data_log_force[1222] <= 18'h1992e;
	 filter_in_data_log_force[1223] <= 18'h1f46e;
	 filter_in_data_log_force[1224] <= 18'h1f373;
	 filter_in_data_log_force[1225] <= 18'h1948d;
	 filter_in_data_log_force[1226] <= 18'h0e7f0;
	 filter_in_data_log_force[1227] <= 18'h00d6d;
	 filter_in_data_log_force[1228] <= 18'h32ee7;
	 filter_in_data_log_force[1229] <= 18'h27876;
	 filter_in_data_log_force[1230] <= 18'h20f92;
	 filter_in_data_log_force[1231] <= 18'h20b1c;
	 filter_in_data_log_force[1232] <= 18'h26df1;
	 filter_in_data_log_force[1233] <= 18'h32560;
	 filter_in_data_log_force[1234] <= 18'h00c2f;
	 filter_in_data_log_force[1235] <= 18'h0f1c4;
	 filter_in_data_log_force[1236] <= 18'h1a43d;
	 filter_in_data_log_force[1237] <= 18'h1fb69;
	 filter_in_data_log_force[1238] <= 18'h1e22d;
	 filter_in_data_log_force[1239] <= 18'h15c2b;
	 filter_in_data_log_force[1240] <= 18'h085f9;
	 filter_in_data_log_force[1241] <= 18'h38f9f;
	 filter_in_data_log_force[1242] <= 18'h2b221;
	 filter_in_data_log_force[1243] <= 18'h2225a;
	 filter_in_data_log_force[1244] <= 18'h2041a;
	 filter_in_data_log_force[1245] <= 18'h260b7;
	 filter_in_data_log_force[1246] <= 18'h323a1;
	 filter_in_data_log_force[1247] <= 18'h01e44;
	 filter_in_data_log_force[1248] <= 18'h112ad;
	 filter_in_data_log_force[1249] <= 18'h1c2af;
	 filter_in_data_log_force[1250] <= 18'h1ffe9;
	 filter_in_data_log_force[1251] <= 18'h1b880;
	 filter_in_data_log_force[1252] <= 18'h0fcfc;
	 filter_in_data_log_force[1253] <= 18'h3fd44;
	 filter_in_data_log_force[1254] <= 18'h2fcf1;
	 filter_in_data_log_force[1255] <= 18'h241af;
	 filter_in_data_log_force[1256] <= 18'h20018;
	 filter_in_data_log_force[1257] <= 18'h24c62;
	 filter_in_data_log_force[1258] <= 18'h3136b;
	 filter_in_data_log_force[1259] <= 18'h01ea4;
	 filter_in_data_log_force[1260] <= 18'h12268;
	 filter_in_data_log_force[1261] <= 18'h1d332;
	 filter_in_data_log_force[1262] <= 18'h1fbd3;
	 filter_in_data_log_force[1263] <= 18'h18e1b;
	 filter_in_data_log_force[1264] <= 18'h0a893;
	 filter_in_data_log_force[1265] <= 18'h38ee2;
	 filter_in_data_log_force[1266] <= 18'h29673;
	 filter_in_data_log_force[1267] <= 18'h20c9e;
	 filter_in_data_log_force[1268] <= 18'h21e24;
	 filter_in_data_log_force[1269] <= 18'h2c7d9;
	 filter_in_data_log_force[1270] <= 18'h3d5e5;
	 filter_in_data_log_force[1271] <= 18'h0f2c3;
	 filter_in_data_log_force[1272] <= 18'h1c1f1;
	 filter_in_data_log_force[1273] <= 18'h1fe28;
	 filter_in_data_log_force[1274] <= 18'h1913e;
	 filter_in_data_log_force[1275] <= 18'h09d42;
	 filter_in_data_log_force[1276] <= 18'h372e9;
	 filter_in_data_log_force[1277] <= 18'h2777d;
	 filter_in_data_log_force[1278] <= 18'h2028d;
	 filter_in_data_log_force[1279] <= 18'h23ed1;
	 filter_in_data_log_force[1280] <= 18'h31994;
	 filter_in_data_log_force[1281] <= 18'h0473f;
	 filter_in_data_log_force[1282] <= 18'h15ca3;
	 filter_in_data_log_force[1283] <= 18'h1f4d3;
	 filter_in_data_log_force[1284] <= 18'h1d65a;
	 filter_in_data_log_force[1285] <= 18'h109f5;
	 filter_in_data_log_force[1286] <= 18'h3d980;
	 filter_in_data_log_force[1287] <= 18'h2b642;
	 filter_in_data_log_force[1288] <= 18'h20f1c;
	 filter_in_data_log_force[1289] <= 18'h225da;
	 filter_in_data_log_force[1290] <= 18'h2f43c;
	 filter_in_data_log_force[1291] <= 18'h02c11;
	 filter_in_data_log_force[1292] <= 18'h153cb;
	 filter_in_data_log_force[1293] <= 18'h1f588;
	 filter_in_data_log_force[1294] <= 18'h1ce94;
	 filter_in_data_log_force[1295] <= 18'h0ec18;
	 filter_in_data_log_force[1296] <= 18'h3a836;
	 filter_in_data_log_force[1297] <= 18'h28742;
	 filter_in_data_log_force[1298] <= 18'h201e8;
	 filter_in_data_log_force[1299] <= 18'h25221;
	 filter_in_data_log_force[1300] <= 18'h358ad;
	 filter_in_data_log_force[1301] <= 18'h0a7b2;
	 filter_in_data_log_force[1302] <= 18'h1afbf;
	 filter_in_data_log_force[1303] <= 18'h1fd2c;
	 filter_in_data_log_force[1304] <= 18'h16bb4;
	 filter_in_data_log_force[1305] <= 18'h038e5;
	 filter_in_data_log_force[1306] <= 18'h2eb93;
	 filter_in_data_log_force[1307] <= 18'h21952;
	 filter_in_data_log_force[1308] <= 18'h222fe;
	 filter_in_data_log_force[1309] <= 18'h306d7;
	 filter_in_data_log_force[1310] <= 18'h05e69;
	 filter_in_data_log_force[1311] <= 18'h18b53;
	 filter_in_data_log_force[1312] <= 18'h1fff8;
	 filter_in_data_log_force[1313] <= 18'h18301;
	 filter_in_data_log_force[1314] <= 18'h04d24;
	 filter_in_data_log_force[1315] <= 18'h2f11e;
	 filter_in_data_log_force[1316] <= 18'h2171a;
	 filter_in_data_log_force[1317] <= 18'h22b18;
	 filter_in_data_log_force[1318] <= 18'h32604;
	 filter_in_data_log_force[1319] <= 18'h08dfc;
	 filter_in_data_log_force[1320] <= 18'h1b027;
	 filter_in_data_log_force[1321] <= 18'h1f965;
	 filter_in_data_log_force[1322] <= 18'h14204;
	 filter_in_data_log_force[1323] <= 18'h3e510;
	 filter_in_data_log_force[1324] <= 18'h294da;
	 filter_in_data_log_force[1325] <= 18'h2007c;
	 filter_in_data_log_force[1326] <= 18'h277dd;
	 filter_in_data_log_force[1327] <= 18'h3bedd;
	 filter_in_data_log_force[1328] <= 18'h1299e;
	 filter_in_data_log_force[1329] <= 18'h1f5d5;
	 filter_in_data_log_force[1330] <= 18'h1b358;
	 filter_in_data_log_force[1331] <= 18'h08370;
	 filter_in_data_log_force[1332] <= 18'h30a67;
	 filter_in_data_log_force[1333] <= 18'h21808;
	 filter_in_data_log_force[1334] <= 18'h234d8;
	 filter_in_data_log_force[1335] <= 18'h3538f;
	 filter_in_data_log_force[1336] <= 18'h0d4b5;
	 filter_in_data_log_force[1337] <= 18'h1ddd4;
	 filter_in_data_log_force[1338] <= 18'h1d574;
	 filter_in_data_log_force[1339] <= 18'h0bd90;
	 filter_in_data_log_force[1340] <= 18'h33665;
	 filter_in_data_log_force[1341] <= 18'h22459;
	 filter_in_data_log_force[1342] <= 18'h22aa0;
	 filter_in_data_log_force[1343] <= 18'h3485b;
	 filter_in_data_log_force[1344] <= 18'h0d50d;
	 filter_in_data_log_force[1345] <= 18'h1e23f;
	 filter_in_data_log_force[1346] <= 18'h1cae8;
	 filter_in_data_log_force[1347] <= 18'h09a62;
	 filter_in_data_log_force[1348] <= 18'h309be;
	 filter_in_data_log_force[1349] <= 18'h210f1;
	 filter_in_data_log_force[1350] <= 18'h24d27;
	 filter_in_data_log_force[1351] <= 18'h39b7e;
	 filter_in_data_log_force[1352] <= 18'h12a89;
	 filter_in_data_log_force[1353] <= 18'h1fbff;
	 filter_in_data_log_force[1354] <= 18'h18749;
	 filter_in_data_log_force[1355] <= 18'h014d8;
	 filter_in_data_log_force[1356] <= 18'h293ca;
	 filter_in_data_log_force[1357] <= 18'h200cc;
	 filter_in_data_log_force[1358] <= 18'h2bf4e;
	 filter_in_data_log_force[1359] <= 18'h053be;
	 filter_in_data_log_force[1360] <= 18'h1b129;
	 filter_in_data_log_force[1361] <= 18'h1eb5e;
	 filter_in_data_log_force[1362] <= 18'h0d81b;
	 filter_in_data_log_force[1363] <= 18'h33069;
	 filter_in_data_log_force[1364] <= 18'h2166f;
	 filter_in_data_log_force[1365] <= 18'h24ec8;
	 filter_in_data_log_force[1366] <= 18'h3b549;
	 filter_in_data_log_force[1367] <= 18'h15123;
	 filter_in_data_log_force[1368] <= 18'h1ffef;
	 filter_in_data_log_force[1369] <= 18'h14340;
	 filter_in_data_log_force[1370] <= 18'h39ecf;
	 filter_in_data_log_force[1371] <= 18'h23f4d;
	 filter_in_data_log_force[1372] <= 18'h22419;
	 filter_in_data_log_force[1373] <= 18'h363f0;
	 filter_in_data_log_force[1374] <= 18'h1171e;
	 filter_in_data_log_force[1375] <= 18'h1fd2f;
	 filter_in_data_log_force[1376] <= 18'h1694e;
	 filter_in_data_log_force[1377] <= 18'h3c6cb;
	 filter_in_data_log_force[1378] <= 18'h24e56;
	 filter_in_data_log_force[1379] <= 18'h21d76;
	 filter_in_data_log_force[1380] <= 18'h35c3f;
	 filter_in_data_log_force[1381] <= 18'h1195e;
	 filter_in_data_log_force[1382] <= 18'h1fe6b;
	 filter_in_data_log_force[1383] <= 18'h157b7;
	 filter_in_data_log_force[1384] <= 18'h3a420;
	 filter_in_data_log_force[1385] <= 18'h237be;
	 filter_in_data_log_force[1386] <= 18'h2334c;
	 filter_in_data_log_force[1387] <= 18'h39d58;
	 filter_in_data_log_force[1388] <= 18'h1572b;
	 filter_in_data_log_force[1389] <= 18'h1fdae;
	 filter_in_data_log_force[1390] <= 18'h107bc;
	 filter_in_data_log_force[1391] <= 18'h33a59;
	 filter_in_data_log_force[1392] <= 18'h20df3;
	 filter_in_data_log_force[1393] <= 18'h27b8f;
	 filter_in_data_log_force[1394] <= 18'h02b94;
	 filter_in_data_log_force[1395] <= 18'h1b82e;
	 filter_in_data_log_force[1396] <= 18'h1d43d;
	 filter_in_data_log_force[1397] <= 18'h06520;
	 filter_in_data_log_force[1398] <= 18'h29f60;
	 filter_in_data_log_force[1399] <= 18'h205c9;
	 filter_in_data_log_force[1400] <= 18'h31ea5;
	 filter_in_data_log_force[1401] <= 18'h0fac1;
	 filter_in_data_log_force[1402] <= 18'h1fe00;
	 filter_in_data_log_force[1403] <= 18'h1442d;
	 filter_in_data_log_force[1404] <= 18'h36d1d;
	 filter_in_data_log_force[1405] <= 18'h216e7;
	 filter_in_data_log_force[1406] <= 18'h272a8;
	 filter_in_data_log_force[1407] <= 18'h031b4;
	 filter_in_data_log_force[1408] <= 18'h1c4f8;
	 filter_in_data_log_force[1409] <= 18'h1bfaa;
	 filter_in_data_log_force[1410] <= 18'h02386;
	 filter_in_data_log_force[1411] <= 18'h2661d;
	 filter_in_data_log_force[1412] <= 18'h2207b;
	 filter_in_data_log_force[1413] <= 18'h395c4;
	 filter_in_data_log_force[1414] <= 18'h16e75;
	 filter_in_data_log_force[1415] <= 18'h1f1bd;
	 filter_in_data_log_force[1416] <= 18'h0a1c9;
	 filter_in_data_log_force[1417] <= 18'h2b86e;
	 filter_in_data_log_force[1418] <= 18'h2052a;
	 filter_in_data_log_force[1419] <= 18'h3355e;
	 filter_in_data_log_force[1420] <= 18'h12898;
	 filter_in_data_log_force[1421] <= 18'h1fe91;
	 filter_in_data_log_force[1422] <= 18'h0e5b1;
	 filter_in_data_log_force[1423] <= 18'h2ec55;
	 filter_in_data_log_force[1424] <= 18'h2004e;
	 filter_in_data_log_force[1425] <= 18'h30c21;
	 filter_in_data_log_force[1426] <= 18'h10a06;
	 filter_in_data_log_force[1427] <= 18'h1ffe2;
	 filter_in_data_log_force[1428] <= 18'h0f5bc;
	 filter_in_data_log_force[1429] <= 18'h2f3d8;
	 filter_in_data_log_force[1430] <= 18'h20052;
	 filter_in_data_log_force[1431] <= 18'h314a2;
	 filter_in_data_log_force[1432] <= 18'h119f6;
	 filter_in_data_log_force[1433] <= 18'h1fe83;
	 filter_in_data_log_force[1434] <= 18'h0d456;
	 filter_in_data_log_force[1435] <= 18'h2cd4f;
	 filter_in_data_log_force[1436] <= 18'h20553;
	 filter_in_data_log_force[1437] <= 18'h35030;
	 filter_in_data_log_force[1438] <= 18'h154d4;
	 filter_in_data_log_force[1439] <= 18'h1f162;
	 filter_in_data_log_force[1440] <= 18'h07cd8;
	 filter_in_data_log_force[1441] <= 18'h28230;
	 filter_in_data_log_force[1442] <= 18'h22125;
	 filter_in_data_log_force[1443] <= 18'h3c53b;
	 filter_in_data_log_force[1444] <= 18'h1a9c4;
	 filter_in_data_log_force[1445] <= 18'h1be90;
	 filter_in_data_log_force[1446] <= 18'h3e9d2;
	 filter_in_data_log_force[1447] <= 18'h22cce;
	 filter_in_data_log_force[1448] <= 18'h27454;
	 filter_in_data_log_force[1449] <= 18'h0741f;
	 filter_in_data_log_force[1450] <= 18'h1f2de;
	 filter_in_data_log_force[1451] <= 18'h141d5;
	 filter_in_data_log_force[1452] <= 18'h3254e;
	 filter_in_data_log_force[1453] <= 18'h20002;
	 filter_in_data_log_force[1454] <= 18'h321b3;
	 filter_in_data_log_force[1455] <= 18'h14252;
	 filter_in_data_log_force[1456] <= 18'h1f0ed;
	 filter_in_data_log_force[1457] <= 18'h0616c;
	 filter_in_data_log_force[1458] <= 18'h2603a;
	 filter_in_data_log_force[1459] <= 18'h2436c;
	 filter_in_data_log_force[1460] <= 18'h02fb7;
	 filter_in_data_log_force[1461] <= 18'h1e47c;
	 filter_in_data_log_force[1462] <= 18'h15c9e;
	 filter_in_data_log_force[1463] <= 18'h3362d;
	 filter_in_data_log_force[1464] <= 18'h20005;
	 filter_in_data_log_force[1465] <= 18'h32faa;
	 filter_in_data_log_force[1466] <= 18'h15acb;
	 filter_in_data_log_force[1467] <= 18'h1e2c5;
	 filter_in_data_log_force[1468] <= 18'h01fc2;
	 filter_in_data_log_force[1469] <= 18'h2355e;
	 filter_in_data_log_force[1470] <= 18'h27d40;
	 filter_in_data_log_force[1471] <= 18'h0a20a;
	 filter_in_data_log_force[1472] <= 18'h1fed5;
	 filter_in_data_log_force[1473] <= 18'h0e094;
	 filter_in_data_log_force[1474] <= 18'h2a959;
	 filter_in_data_log_force[1475] <= 18'h21f83;
	 filter_in_data_log_force[1476] <= 18'h3f348;
	 filter_in_data_log_force[1477] <= 18'h1d7b7;
	 filter_in_data_log_force[1478] <= 18'h164bb;
	 filter_in_data_log_force[1479] <= 18'h329e1;
	 filter_in_data_log_force[1480] <= 18'h2011d;
	 filter_in_data_log_force[1481] <= 18'h36a6c;
	 filter_in_data_log_force[1482] <= 18'h195c0;
	 filter_in_data_log_force[1483] <= 18'h1b239;
	 filter_in_data_log_force[1484] <= 18'h397c8;
	 filter_in_data_log_force[1485] <= 18'h20568;
	 filter_in_data_log_force[1486] <= 18'h30dc0;
	 filter_in_data_log_force[1487] <= 18'h156c8;
	 filter_in_data_log_force[1488] <= 18'h1d923;
	 filter_in_data_log_force[1489] <= 18'h3e47f;
	 filter_in_data_log_force[1490] <= 18'h2142c;
	 filter_in_data_log_force[1491] <= 18'h2d903;
	 filter_in_data_log_force[1492] <= 18'h12c94;
	 filter_in_data_log_force[1493] <= 18'h1e8f8;
	 filter_in_data_log_force[1494] <= 18'h00b66;
	 filter_in_data_log_force[1495] <= 18'h21dc1;
	 filter_in_data_log_force[1496] <= 18'h2c61e;
	 filter_in_data_log_force[1497] <= 18'h11fa5;
	 filter_in_data_log_force[1498] <= 18'h1eb4f;
	 filter_in_data_log_force[1499] <= 18'h00bcb;
	 filter_in_data_log_force[1500] <= 18'h21b59;
	 filter_in_data_log_force[1501] <= 18'h2d21d;
	 filter_in_data_log_force[1502] <= 18'h13226;
	 filter_in_data_log_force[1503] <= 18'h1e1e3;
	 filter_in_data_log_force[1504] <= 18'h3e5ad;
	 filter_in_data_log_force[1505] <= 18'h20e87;
	 filter_in_data_log_force[1506] <= 18'h2feed;
	 filter_in_data_log_force[1507] <= 18'h160ef;
	 filter_in_data_log_force[1508] <= 18'h1c64c;
	 filter_in_data_log_force[1509] <= 18'h399b5;
	 filter_in_data_log_force[1510] <= 18'h20167;
	 filter_in_data_log_force[1511] <= 18'h35241;
	 filter_in_data_log_force[1512] <= 18'h1a213;
	 filter_in_data_log_force[1513] <= 18'h18b20;
	 filter_in_data_log_force[1514] <= 18'h32c61;
	 filter_in_data_log_force[1515] <= 18'h20709;
	 filter_in_data_log_force[1516] <= 18'h3d162;
	 filter_in_data_log_force[1517] <= 18'h1e1c7;
	 filter_in_data_log_force[1518] <= 18'h11f94;
	 filter_in_data_log_force[1519] <= 18'h2abfc;
	 filter_in_data_log_force[1520] <= 18'h23a24;
	 filter_in_data_log_force[1521] <= 18'h07942;
	 filter_in_data_log_force[1522] <= 18'h1ffff;
	 filter_in_data_log_force[1523] <= 18'h077bb;
	 filter_in_data_log_force[1524] <= 18'h2374e;
	 filter_in_data_log_force[1525] <= 18'h2b680;
	 filter_in_data_log_force[1526] <= 18'h133a9;
	 filter_in_data_log_force[1527] <= 18'h1d360;
	 filter_in_data_log_force[1528] <= 18'h39a7e;
	 filter_in_data_log_force[1529] <= 18'h20016;
	 filter_in_data_log_force[1530] <= 18'h38992;
	 filter_in_data_log_force[1531] <= 18'h1ce0c;
	 filter_in_data_log_force[1532] <= 18'h137a4;
	 filter_in_data_log_force[1533] <= 18'h2b218;
	 filter_in_data_log_force[1534] <= 18'h24087;
	 filter_in_data_log_force[1535] <= 18'h09afc;
	 filter_in_data_log_force[1536] <= 18'h1fcdf;
	 filter_in_data_log_force[1537] <= 18'h02aa0;
	 filter_in_data_log_force[1538] <= 18'h21323;
	 filter_in_data_log_force[1539] <= 18'h31bb3;
	 filter_in_data_log_force[1540] <= 18'h1987f;
	 filter_in_data_log_force[1541] <= 18'h17977;
	 filter_in_data_log_force[1542] <= 18'h2eec2;
	 filter_in_data_log_force[1543] <= 18'h225e1;
	 filter_in_data_log_force[1544] <= 18'h06cd5;
	 filter_in_data_log_force[1545] <= 18'h1ff7f;
	 filter_in_data_log_force[1546] <= 18'h03e90;
	 filter_in_data_log_force[1547] <= 18'h214d9;
	 filter_in_data_log_force[1548] <= 18'h3229b;
	 filter_in_data_log_force[1549] <= 18'h1a521;
	 filter_in_data_log_force[1550] <= 18'h160a6;
	 filter_in_data_log_force[1551] <= 18'h2c667;
	 filter_in_data_log_force[1552] <= 18'h24143;
	 filter_in_data_log_force[1553] <= 18'h0b697;
	 filter_in_data_log_force[1554] <= 18'h1f373;
	 filter_in_data_log_force[1555] <= 18'h3d601;
	 filter_in_data_log_force[1556] <= 18'h200c4;
	 filter_in_data_log_force[1557] <= 18'h3a01f;
	 filter_in_data_log_force[1558] <= 18'h1e627;
	 filter_in_data_log_force[1559] <= 18'h0dd3d;
	 filter_in_data_log_force[1560] <= 18'h2515f;
	 filter_in_data_log_force[1561] <= 18'h2b8d1;
	 filter_in_data_log_force[1562] <= 18'h1604e;
	 filter_in_data_log_force[1563] <= 18'h199b3;
	 filter_in_data_log_force[1564] <= 18'h2fcf1;
	 filter_in_data_log_force[1565] <= 18'h22cad;
	 filter_in_data_log_force[1566] <= 18'h09e3b;
	 filter_in_data_log_force[1567] <= 18'h1f4b2;
	 filter_in_data_log_force[1568] <= 18'h3c7d7;
	 filter_in_data_log_force[1569] <= 18'h2000a;
	 filter_in_data_log_force[1570] <= 18'h3d5e5;
	 filter_in_data_log_force[1571] <= 18'h1f846;
	 filter_in_data_log_force[1572] <= 18'h084e1;
	 filter_in_data_log_force[1573] <= 18'h21eb6;
	 filter_in_data_log_force[1574] <= 18'h32a3c;
	 filter_in_data_log_force[1575] <= 18'h1bec7;
	 filter_in_data_log_force[1576] <= 18'h11b82;
	 filter_in_data_log_force[1577] <= 18'h26ba5;
	 filter_in_data_log_force[1578] <= 18'h2aa36;
	 filter_in_data_log_force[1579] <= 18'h16548;
	 filter_in_data_log_force[1580] <= 18'h18502;
	 filter_in_data_log_force[1581] <= 18'h2cba6;
	 filter_in_data_log_force[1582] <= 18'h255f0;
	 filter_in_data_log_force[1583] <= 18'h103db;
	 filter_in_data_log_force[1584] <= 18'h1c62e;
	 filter_in_data_log_force[1585] <= 18'h32a64;
	 filter_in_data_log_force[1586] <= 18'h22545;
	 filter_in_data_log_force[1587] <= 18'h0aaf6;
	 filter_in_data_log_force[1588] <= 18'h1e922;
	 filter_in_data_log_force[1589] <= 18'h37b1b;
	 filter_in_data_log_force[1590] <= 18'h20d44;
	 filter_in_data_log_force[1591] <= 18'h06413;
	 filter_in_data_log_force[1592] <= 18'h1f8c4;
	 filter_in_data_log_force[1593] <= 18'h3b713;
	 filter_in_data_log_force[1594] <= 18'h203b7;
	 filter_in_data_log_force[1595] <= 18'h033b4;
	 filter_in_data_log_force[1596] <= 18'h1fe29;
	 filter_in_data_log_force[1597] <= 18'h3db75;
	 filter_in_data_log_force[1598] <= 18'h200f4;
	 filter_in_data_log_force[1599] <= 18'h01b81;
	 filter_in_data_log_force[1600] <= 18'h1ff60;
	 filter_in_data_log_force[1601] <= 18'h3e763;
	 filter_in_data_log_force[1602] <= 18'h200a2;
	 filter_in_data_log_force[1603] <= 18'h01be1;
	 filter_in_data_log_force[1604] <= 18'h1ff03;
	 filter_in_data_log_force[1605] <= 18'h3dab5;
	 filter_in_data_log_force[1606] <= 18'h201ec;
	 filter_in_data_log_force[1607] <= 18'h034d5;
	 filter_in_data_log_force[1608] <= 18'h1fc20;
	 filter_in_data_log_force[1609] <= 18'h3b594;
	 filter_in_data_log_force[1610] <= 18'h20786;
	 filter_in_data_log_force[1611] <= 18'h065ed;
	 filter_in_data_log_force[1612] <= 18'h1f242;
	 filter_in_data_log_force[1613] <= 18'h378eb;
	 filter_in_data_log_force[1614] <= 18'h21799;
	 filter_in_data_log_force[1615] <= 18'h0ad73;
	 filter_in_data_log_force[1616] <= 18'h1d9aa;
	 filter_in_data_log_force[1617] <= 18'h327a7;
	 filter_in_data_log_force[1618] <= 18'h23b4f;
	 filter_in_data_log_force[1619] <= 18'h106c7;
	 filter_in_data_log_force[1620] <= 18'h1a811;
	 filter_in_data_log_force[1621] <= 18'h2c8a5;
	 filter_in_data_log_force[1622] <= 18'h27d95;
	 filter_in_data_log_force[1623] <= 18'h1683f;
	 filter_in_data_log_force[1624] <= 18'h1528b;
	 filter_in_data_log_force[1625] <= 18'h268e2;
	 filter_in_data_log_force[1626] <= 18'h2e86f;
	 filter_in_data_log_force[1627] <= 18'h1c127;
	 filter_in_data_log_force[1628] <= 18'h0d120;
	 filter_in_data_log_force[1629] <= 18'h21cf0;
	 filter_in_data_log_force[1630] <= 18'h38069;
	 filter_in_data_log_force[1631] <= 18'h1f939;
	 filter_in_data_log_force[1632] <= 18'h02446;
	 filter_in_data_log_force[1633] <= 18'h20026;
	 filter_in_data_log_force[1634] <= 18'h03e58;
	 filter_in_data_log_force[1635] <= 18'h1f350;
	 filter_in_data_log_force[1636] <= 18'h35b80;
	 filter_in_data_log_force[1637] <= 18'h22f7e;
	 filter_in_data_log_force[1638] <= 18'h1090e;
	 filter_in_data_log_force[1639] <= 18'h1955c;
	 filter_in_data_log_force[1640] <= 18'h29a64;
	 filter_in_data_log_force[1641] <= 18'h2bea8;
	 filter_in_data_log_force[1642] <= 18'h1b2c3;
	 filter_in_data_log_force[1643] <= 18'h0d611;
	 filter_in_data_log_force[1644] <= 18'h2175d;
	 filter_in_data_log_force[1645] <= 18'h3a84a;
	 filter_in_data_log_force[1646] <= 18'h1ffa1;
	 filter_in_data_log_force[1647] <= 18'h3cd5c;
	 filter_in_data_log_force[1648] <= 18'h20e94;
	 filter_in_data_log_force[1649] <= 18'h0bf05;
	 filter_in_data_log_force[1650] <= 18'h1ba26;
	 filter_in_data_log_force[1651] <= 18'h2bf00;
	 filter_in_data_log_force[1652] <= 18'h2a664;
	 filter_in_data_log_force[1653] <= 18'h1aaa1;
	 filter_in_data_log_force[1654] <= 18'h0d456;
	 filter_in_data_log_force[1655] <= 18'h21211;
	 filter_in_data_log_force[1656] <= 18'h3cbc0;
	 filter_in_data_log_force[1657] <= 18'h1feeb;
	 filter_in_data_log_force[1658] <= 18'h388af;
	 filter_in_data_log_force[1659] <= 18'h22a1e;
	 filter_in_data_log_force[1660] <= 18'h11a97;
	 filter_in_data_log_force[1661] <= 18'h171ba;
	 filter_in_data_log_force[1662] <= 18'h260ab;
	 filter_in_data_log_force[1663] <= 18'h3263b;
	 filter_in_data_log_force[1664] <= 18'h1eff3;
	 filter_in_data_log_force[1665] <= 18'h01e94;
	 filter_in_data_log_force[1666] <= 18'h204a0;
	 filter_in_data_log_force[1667] <= 18'h0a6ce;
	 filter_in_data_log_force[1668] <= 18'h1b932;
	 filter_in_data_log_force[1669] <= 18'h2a879;
	 filter_in_data_log_force[1670] <= 18'h2d2c9;
	 filter_in_data_log_force[1671] <= 18'h1d395;
	 filter_in_data_log_force[1672] <= 18'h0695c;
	 filter_in_data_log_force[1673] <= 18'h20004;
	 filter_in_data_log_force[1674] <= 18'h072f8;
	 filter_in_data_log_force[1675] <= 18'h1cd81;
	 filter_in_data_log_force[1676] <= 18'h2c126;
	 filter_in_data_log_force[1677] <= 18'h2c19a;
	 filter_in_data_log_force[1678] <= 18'h1cf14;
	 filter_in_data_log_force[1679] <= 18'h06960;
	 filter_in_data_log_force[1680] <= 18'h20038;
	 filter_in_data_log_force[1681] <= 18'h087de;
	 filter_in_data_log_force[1682] <= 18'h1be96;
	 filter_in_data_log_force[1683] <= 18'h2a093;
	 filter_in_data_log_force[1684] <= 18'h2ed83;
	 filter_in_data_log_force[1685] <= 18'h1e6e9;
	 filter_in_data_log_force[1686] <= 18'h01ea0;
	 filter_in_data_log_force[1687] <= 18'h209f8;
	 filter_in_data_log_force[1688] <= 18'h0e275;
	 filter_in_data_log_force[1689] <= 18'h1805c;
	 filter_in_data_log_force[1690] <= 18'h25476;
	 filter_in_data_log_force[1691] <= 18'h36252;
	 filter_in_data_log_force[1692] <= 18'h1ff94;
	 filter_in_data_log_force[1693] <= 18'h388c2;
	 filter_in_data_log_force[1694] <= 18'h24210;
	 filter_in_data_log_force[1695] <= 18'h16d91;
	 filter_in_data_log_force[1696] <= 18'h0f16b;
	 filter_in_data_log_force[1697] <= 18'h20a8f;
	 filter_in_data_log_force[1698] <= 18'h02c95;
	 filter_in_data_log_force[1699] <= 18'h1db53;
	 filter_in_data_log_force[1700] <= 18'h2bf16;
	 filter_in_data_log_force[1701] <= 18'h2e18e;
	 filter_in_data_log_force[1702] <= 18'h1ea76;
	 filter_in_data_log_force[1703] <= 18'h3f88c;
	 filter_in_data_log_force[1704] <= 18'h21a83;
	 filter_in_data_log_force[1705] <= 18'h12fa9;
	 filter_in_data_log_force[1706] <= 18'h12a00;
	 filter_in_data_log_force[1707] <= 18'h21768;
	 filter_in_data_log_force[1708] <= 18'h008ca;
	 filter_in_data_log_force[1709] <= 18'h1e28a;
	 filter_in_data_log_force[1710] <= 18'h2c305;
	 filter_in_data_log_force[1711] <= 18'h2ea37;
	 filter_in_data_log_force[1712] <= 18'h1f13c;
	 filter_in_data_log_force[1713] <= 18'h3cf6d;
	 filter_in_data_log_force[1714] <= 18'h22f6b;
	 filter_in_data_log_force[1715] <= 18'h16674;
	 filter_in_data_log_force[1716] <= 18'h0deec;
	 filter_in_data_log_force[1717] <= 18'h202b3;
	 filter_in_data_log_force[1718] <= 18'h07dbb;
	 filter_in_data_log_force[1719] <= 18'h1a605;
	 filter_in_data_log_force[1720] <= 18'h25cf3;
	 filter_in_data_log_force[1721] <= 18'h38037;
	 filter_in_data_log_force[1722] <= 18'h1fcdf;
	 filter_in_data_log_force[1723] <= 18'h31531;
	 filter_in_data_log_force[1724] <= 18'h2ac47;
	 filter_in_data_log_force[1725] <= 18'h1e051;
	 filter_in_data_log_force[1726] <= 18'h3f523;
	 filter_in_data_log_force[1727] <= 18'h2283d;
	 filter_in_data_log_force[1728] <= 18'h16814;
	 filter_in_data_log_force[1729] <= 18'h0caa2;
	 filter_in_data_log_force[1730] <= 18'h2001a;
	 filter_in_data_log_force[1731] <= 18'h0b91d;
	 filter_in_data_log_force[1732] <= 18'h1721b;
	 filter_in_data_log_force[1733] <= 18'h22ad8;
	 filter_in_data_log_force[1734] <= 18'h3f951;
	 filter_in_data_log_force[1735] <= 18'h1d9c4;
	 filter_in_data_log_force[1736] <= 18'h292e8;
	 filter_in_data_log_force[1737] <= 18'h3475b;
	 filter_in_data_log_force[1738] <= 18'h1ff8c;
	 filter_in_data_log_force[1739] <= 18'h31e85;
	 filter_in_data_log_force[1740] <= 18'h2b70b;
	 filter_in_data_log_force[1741] <= 18'h1ec61;
	 filter_in_data_log_force[1742] <= 18'h3b5e0;
	 filter_in_data_log_force[1743] <= 18'h25150;
	 filter_in_data_log_force[1744] <= 18'h1aeef;
	 filter_in_data_log_force[1745] <= 18'h046a0;
	 filter_in_data_log_force[1746] <= 18'h2165e;
	 filter_in_data_log_force[1747] <= 18'h15740;
	 filter_in_data_log_force[1748] <= 18'h0c500;
	 filter_in_data_log_force[1749] <= 18'h2009e;
	 filter_in_data_log_force[1750] <= 18'h0f3c6;
	 filter_in_data_log_force[1751] <= 18'h12b57;
	 filter_in_data_log_force[1752] <= 18'h2077f;
	 filter_in_data_log_force[1753] <= 18'h08fdb;
	 filter_in_data_log_force[1754] <= 18'h178bc;
	 filter_in_data_log_force[1755] <= 18'h221ad;
	 filter_in_data_log_force[1756] <= 18'h03358;
	 filter_in_data_log_force[1757] <= 18'h1af6f;
	 filter_in_data_log_force[1758] <= 18'h24680;
	 filter_in_data_log_force[1759] <= 18'h3e2ed;
	 filter_in_data_log_force[1760] <= 18'h1d36c;
	 filter_in_data_log_force[1761] <= 18'h26ec0;
	 filter_in_data_log_force[1762] <= 18'h3a0d1;
	 filter_in_data_log_force[1763] <= 18'h1e93f;
	 filter_in_data_log_force[1764] <= 18'h294da;
	 filter_in_data_log_force[1765] <= 18'h36d8d;
	 filter_in_data_log_force[1766] <= 18'h1f543;
	 filter_in_data_log_force[1767] <= 18'h2b4d1;
	 filter_in_data_log_force[1768] <= 18'h348b9;
	 filter_in_data_log_force[1769] <= 18'h1fb1e;
	 filter_in_data_log_force[1770] <= 18'h2cbfd;
	 filter_in_data_log_force[1771] <= 18'h33190;
	 filter_in_data_log_force[1772] <= 18'h1fd87;
	 filter_in_data_log_force[1773] <= 18'h2d8c1;
	 filter_in_data_log_force[1774] <= 18'h32762;
	 filter_in_data_log_force[1775] <= 18'h1fe21;
	 filter_in_data_log_force[1776] <= 18'h2da56;
	 filter_in_data_log_force[1777] <= 18'h329d2;
	 filter_in_data_log_force[1778] <= 18'h1fd74;
	 filter_in_data_log_force[1779] <= 18'h2d0a4;
	 filter_in_data_log_force[1780] <= 18'h338f8;
	 filter_in_data_log_force[1781] <= 18'h1fae9;
	 filter_in_data_log_force[1782] <= 18'h2bc40;
	 filter_in_data_log_force[1783] <= 18'h35556;
	 filter_in_data_log_force[1784] <= 18'h1f4cc;
	 filter_in_data_log_force[1785] <= 18'h29e85;
	 filter_in_data_log_force[1786] <= 18'h37fae;
	 filter_in_data_log_force[1787] <= 18'h1e859;
	 filter_in_data_log_force[1788] <= 18'h279ca;
	 filter_in_data_log_force[1789] <= 18'h3b8b1;
	 filter_in_data_log_force[1790] <= 18'h1d1de;
	 filter_in_data_log_force[1791] <= 18'h251a7;
	 filter_in_data_log_force[1792] <= 18'h0007d;
	 filter_in_data_log_force[1793] <= 18'h1acfb;
	 filter_in_data_log_force[1794] <= 18'h22b37;
	 filter_in_data_log_force[1795] <= 18'h055fa;
	 filter_in_data_log_force[1796] <= 18'h17523;
	 filter_in_data_log_force[1797] <= 18'h20d40;
	 filter_in_data_log_force[1798] <= 18'h0b613;
	 filter_in_data_log_force[1799] <= 18'h1266c;
	 filter_in_data_log_force[1800] <= 18'h2000f;
	 filter_in_data_log_force[1801] <= 18'h11af2;
	 filter_in_data_log_force[1802] <= 18'h0beb7;
	 filter_in_data_log_force[1803] <= 18'h20ce5;
	 filter_in_data_log_force[1804] <= 18'h17b62;
	 filter_in_data_log_force[1805] <= 18'h03f24;
	 filter_in_data_log_force[1806] <= 18'h23cba;
	 filter_in_data_log_force[1807] <= 18'h1cabf;
	 filter_in_data_log_force[1808] <= 18'h3adac;
	 filter_in_data_log_force[1809] <= 18'h2963d;
	 filter_in_data_log_force[1810] <= 18'h1f9b5;
	 filter_in_data_log_force[1811] <= 18'h3166c;
	 filter_in_data_log_force[1812] <= 18'h31b27;
	 filter_in_data_log_force[1813] <= 18'h1f854;
	 filter_in_data_log_force[1814] <= 18'h28c18;
	 filter_in_data_log_force[1815] <= 18'h3c53b;
	 filter_in_data_log_force[1816] <= 18'h1b994;
	 filter_in_data_log_force[1817] <= 18'h226b6;
	 filter_in_data_log_force[1818] <= 18'h083d1;
	 filter_in_data_log_force[1819] <= 18'h13827;
	 filter_in_data_log_force[1820] <= 18'h20000;
	 filter_in_data_log_force[1821] <= 18'h13b16;
	 filter_in_data_log_force[1822] <= 18'h07bbf;
	 filter_in_data_log_force[1823] <= 18'h22d10;
	 filter_in_data_log_force[1824] <= 18'h1c68b;
	 filter_in_data_log_force[1825] <= 18'h39d09;
	 filter_in_data_log_force[1826] <= 18'h2b5fb;
	 filter_in_data_log_force[1827] <= 18'h1ffe1;
	 filter_in_data_log_force[1828] <= 18'h2c5fe;
	 filter_in_data_log_force[1829] <= 18'h38d6a;
	 filter_in_data_log_force[1830] <= 18'h1ca4a;
	 filter_in_data_log_force[1831] <= 18'h22c09;
	 filter_in_data_log_force[1832] <= 18'h08b94;
	 filter_in_data_log_force[1833] <= 18'h1202a;
	 filter_in_data_log_force[1834] <= 18'h202ab;
	 filter_in_data_log_force[1835] <= 18'h17113;
	 filter_in_data_log_force[1836] <= 18'h01ea0;
	 filter_in_data_log_force[1837] <= 18'h2681f;
	 filter_in_data_log_force[1838] <= 18'h1f4c7;
	 filter_in_data_log_force[1839] <= 18'h30837;
	 filter_in_data_log_force[1840] <= 18'h35190;
	 filter_in_data_log_force[1841] <= 18'h1dcbd;
	 filter_in_data_log_force[1842] <= 18'h23856;
	 filter_in_data_log_force[1843] <= 18'h08065;
	 filter_in_data_log_force[1844] <= 18'h11bb7;
	 filter_in_data_log_force[1845] <= 18'h2056d;
	 filter_in_data_log_force[1846] <= 18'h18b2c;
	 filter_in_data_log_force[1847] <= 18'h3e672;
	 filter_in_data_log_force[1848] <= 18'h29859;
	 filter_in_data_log_force[1849] <= 18'h1ffb5;
	 filter_in_data_log_force[1850] <= 18'h2b09b;
	 filter_in_data_log_force[1851] <= 18'h3ca1b;
	 filter_in_data_log_force[1852] <= 18'h19806;
	 filter_in_data_log_force[1853] <= 18'h206f6;
	 filter_in_data_log_force[1854] <= 18'h11efb;
	 filter_in_data_log_force[1855] <= 18'h06c15;
	 filter_in_data_log_force[1856] <= 18'h24c6d;
	 filter_in_data_log_force[1857] <= 18'h1f04e;
	 filter_in_data_log_force[1858] <= 18'h2ffe1;
	 filter_in_data_log_force[1859] <= 18'h3768e;
	 filter_in_data_log_force[1860] <= 18'h1bfc0;
	 filter_in_data_log_force[1861] <= 18'h21467;
	 filter_in_data_log_force[1862] <= 18'h0f5df;
	 filter_in_data_log_force[1863] <= 18'h08ed4;
	 filter_in_data_log_force[1864] <= 18'h24087;
	 filter_in_data_log_force[1865] <= 18'h1ed6f;
	 filter_in_data_log_force[1866] <= 18'h2fee6;
	 filter_in_data_log_force[1867] <= 18'h38391;
	 filter_in_data_log_force[1868] <= 18'h1b2ae;
	 filter_in_data_log_force[1869] <= 18'h20b20;
	 filter_in_data_log_force[1870] <= 18'h120da;
	 filter_in_data_log_force[1871] <= 18'h051a2;
	 filter_in_data_log_force[1872] <= 18'h269b1;
	 filter_in_data_log_force[1873] <= 18'h1fd79;
	 filter_in_data_log_force[1874] <= 18'h2ae0c;
	 filter_in_data_log_force[1875] <= 18'h3f263;
	 filter_in_data_log_force[1876] <= 18'h164d2;
	 filter_in_data_log_force[1877] <= 18'h200de;
	 filter_in_data_log_force[1878] <= 18'h18e0a;
	 filter_in_data_log_force[1879] <= 18'h3b0ea;
	 filter_in_data_log_force[1880] <= 18'h2e88a;
	 filter_in_data_log_force[1881] <= 18'h1ee44;
	 filter_in_data_log_force[1882] <= 18'h235c8;
	 filter_in_data_log_force[1883] <= 18'h0c03f;
	 filter_in_data_log_force[1884] <= 18'h0a893;
	 filter_in_data_log_force[1885] <= 18'h24324;
	 filter_in_data_log_force[1886] <= 18'h1f625;
	 filter_in_data_log_force[1887] <= 18'h2c4ea;
	 filter_in_data_log_force[1888] <= 18'h3e8b9;
	 filter_in_data_log_force[1889] <= 18'h15d51;
	 filter_in_data_log_force[1890] <= 18'h20389;
	 filter_in_data_log_force[1891] <= 18'h1abc6;
	 filter_in_data_log_force[1892] <= 18'h36c46;
	 filter_in_data_log_force[1893] <= 18'h33851;
	 filter_in_data_log_force[1894] <= 18'h1c62e;
	 filter_in_data_log_force[1895] <= 18'h20afb;
	 filter_in_data_log_force[1896] <= 18'h1418d;
	 filter_in_data_log_force[1897] <= 18'h0012a;
	 filter_in_data_log_force[1898] <= 18'h2bdd6;
	 filter_in_data_log_force[1899] <= 18'h1f437;
	 filter_in_data_log_force[1900] <= 18'h2349c;
	 filter_in_data_log_force[1901] <= 18'h0dc0c;
	 filter_in_data_log_force[1902] <= 18'h070bc;
	 filter_in_data_log_force[1903] <= 18'h273ae;
	 filter_in_data_log_force[1904] <= 18'h1ffd6;
	 filter_in_data_log_force[1905] <= 18'h262dc;
	 filter_in_data_log_force[1906] <= 18'h08fcf;
	 filter_in_data_log_force[1907] <= 18'h0b778;
	 filter_in_data_log_force[1908] <= 18'h24d27;
	 filter_in_data_log_force[1909] <= 18'h1fdf9;
	 filter_in_data_log_force[1910] <= 18'h282e4;
	 filter_in_data_log_force[1911] <= 18'h065ed;
	 filter_in_data_log_force[1912] <= 18'h0d81b;
	 filter_in_data_log_force[1913] <= 18'h23f26;
	 filter_in_data_log_force[1914] <= 18'h1fbcc;
	 filter_in_data_log_force[1915] <= 18'h28b3e;
	 filter_in_data_log_force[1916] <= 18'h06160;
	 filter_in_data_log_force[1917] <= 18'h0d552;
	 filter_in_data_log_force[1918] <= 18'h2446e;
	 filter_in_data_log_force[1919] <= 18'h1fdd4;
	 filter_in_data_log_force[1920] <= 18'h279ca;
	 filter_in_data_log_force[1921] <= 18'h08267;
	 filter_in_data_log_force[1922] <= 18'h0aeda;
	 filter_in_data_log_force[1923] <= 18'h25f11;
	 filter_in_data_log_force[1924] <= 18'h1ffe8;
	 filter_in_data_log_force[1925] <= 18'h25320;
	 filter_in_data_log_force[1926] <= 18'h0c6e3;
	 filter_in_data_log_force[1927] <= 18'h061bb;
	 filter_in_data_log_force[1928] <= 18'h297e7;
	 filter_in_data_log_force[1929] <= 18'h1f533;
	 filter_in_data_log_force[1930] <= 18'h223cf;
	 filter_in_data_log_force[1931] <= 18'h127a8;
	 filter_in_data_log_force[1932] <= 18'h3ebb5;
	 filter_in_data_log_force[1933] <= 18'h2fbb6;
	 filter_in_data_log_force[1934] <= 18'h1c90d;
	 filter_in_data_log_force[1935] <= 18'h20287;
	 filter_in_data_log_force[1936] <= 18'h19370;
	 filter_in_data_log_force[1937] <= 18'h35214;
	 filter_in_data_log_force[1938] <= 18'h3949c;
	 filter_in_data_log_force[1939] <= 18'h16306;
	 filter_in_data_log_force[1940] <= 18'h21043;
	 filter_in_data_log_force[1941] <= 18'h1e9b6;
	 filter_in_data_log_force[1942] <= 18'h2ab08;
	 filter_in_data_log_force[1943] <= 18'h05ea4;
	 filter_in_data_log_force[1944] <= 18'h0b174;
	 filter_in_data_log_force[1945] <= 18'h271e5;
	 filter_in_data_log_force[1946] <= 18'h1fa8a;
	 filter_in_data_log_force[1947] <= 18'h22567;
	 filter_in_data_log_force[1948] <= 18'h13943;
	 filter_in_data_log_force[1949] <= 18'h3bbcf;
	 filter_in_data_log_force[1950] <= 18'h33e32;
	 filter_in_data_log_force[1951] <= 18'h19346;
	 filter_in_data_log_force[1952] <= 18'h2059a;
	 filter_in_data_log_force[1953] <= 18'h1de53;
	 filter_in_data_log_force[1954] <= 18'h2b799;
	 filter_in_data_log_force[1955] <= 18'h0607f;
	 filter_in_data_log_force[1956] <= 18'h09e34;
	 filter_in_data_log_force[1957] <= 18'h28b75;
	 filter_in_data_log_force[1958] <= 18'h1ef06;
	 filter_in_data_log_force[1959] <= 18'h20e3f;
	 filter_in_data_log_force[1960] <= 18'h17e29;
	 filter_in_data_log_force[1961] <= 18'h34e89;
	 filter_in_data_log_force[1962] <= 18'h3bcc2;
	 filter_in_data_log_force[1963] <= 18'h12724;
	 filter_in_data_log_force[1964] <= 18'h23919;
	 filter_in_data_log_force[1965] <= 18'h1ffff;
	 filter_in_data_log_force[1966] <= 18'h23856;
	 filter_in_data_log_force[1967] <= 18'h12c42;
	 filter_in_data_log_force[1968] <= 18'h3aee9;
	 filter_in_data_log_force[1969] <= 18'h365fa;
	 filter_in_data_log_force[1970] <= 18'h16360;
	 filter_in_data_log_force[1971] <= 18'h21e2e;
	 filter_in_data_log_force[1972] <= 18'h1fce0;
	 filter_in_data_log_force[1973] <= 18'h24f0c;
	 filter_in_data_log_force[1974] <= 18'h10f2a;
	 filter_in_data_log_force[1975] <= 18'h3c6fb;
	 filter_in_data_log_force[1976] <= 18'h35927;
	 filter_in_data_log_force[1977] <= 18'h16554;
	 filter_in_data_log_force[1978] <= 18'h220f7;
	 filter_in_data_log_force[1979] <= 18'h1fe9c;
	 filter_in_data_log_force[1980] <= 18'h23ff6;
	 filter_in_data_log_force[1981] <= 18'h13093;
	 filter_in_data_log_force[1982] <= 18'h39475;
	 filter_in_data_log_force[1983] <= 18'h394d8;
	 filter_in_data_log_force[1984] <= 18'h12dc6;
	 filter_in_data_log_force[1985] <= 18'h244b5;
	 filter_in_data_log_force[1986] <= 18'h1fcdf;
	 filter_in_data_log_force[1987] <= 18'h216d8;
	 filter_in_data_log_force[1988] <= 18'h18531;
	 filter_in_data_log_force[1989] <= 18'h31d1c;
	 filter_in_data_log_force[1990] <= 18'h01d87;
	 filter_in_data_log_force[1991] <= 18'h0ab14;
	 filter_in_data_log_force[1992] <= 18'h2a840;
	 filter_in_data_log_force[1993] <= 18'h1ceb9;
	 filter_in_data_log_force[1994] <= 18'h200b8;
	 filter_in_data_log_force[1995] <= 18'h1e3cf;
	 filter_in_data_log_force[1996] <= 18'h27df9;
	 filter_in_data_log_force[1997] <= 18'h0e994;
	 filter_in_data_log_force[1998] <= 18'h3ceb9;
	 filter_in_data_log_force[1999] <= 18'h37387;
	 filter_in_data_log_force[2000] <= 18'h1358b;
	 filter_in_data_log_force[2001] <= 18'h24c62;
	 filter_in_data_log_force[2002] <= 18'h1f6fb;
	 filter_in_data_log_force[2003] <= 18'h207c2;
	 filter_in_data_log_force[2004] <= 18'h1b8d4;
	 filter_in_data_log_force[2005] <= 18'h2bdae;
	 filter_in_data_log_force[2006] <= 18'h0a4cc;
	 filter_in_data_log_force[2007] <= 18'h00b8a;
	 filter_in_data_log_force[2008] <= 18'h346f6;
	 filter_in_data_log_force[2009] <= 18'h14f4a;
	 filter_in_data_log_force[2010] <= 18'h2428f;
	 filter_in_data_log_force[2011] <= 18'h1f7f7;
	 filter_in_data_log_force[2012] <= 18'h2065d;
	 filter_in_data_log_force[2013] <= 18'h1c3c1;
	 filter_in_data_log_force[2014] <= 18'h2a265;
	 filter_in_data_log_force[2015] <= 18'h0d352;
	 filter_in_data_log_force[2016] <= 18'h3cbb8;
	 filter_in_data_log_force[2017] <= 18'h39157;
	 filter_in_data_log_force[2018] <= 18'h10509;
	 filter_in_data_log_force[2019] <= 18'h27fa4;
	 filter_in_data_log_force[2020] <= 18'h1d574;
	 filter_in_data_log_force[2021] <= 18'h202af;
	 filter_in_data_log_force[2022] <= 18'h1f586;
	 filter_in_data_log_force[2023] <= 18'h23fd9;
	 filter_in_data_log_force[2024] <= 18'h1634f;
	 filter_in_data_log_force[2025] <= 18'h317b6;
	 filter_in_data_log_force[2026] <= 18'h05a93;
	 filter_in_data_log_force[2027] <= 18'h03955;
	 filter_in_data_log_force[2028] <= 18'h338f8;
	 filter_in_data_log_force[2029] <= 18'h14340;
	 filter_in_data_log_force[2030] <= 18'h25b50;
	 filter_in_data_log_force[2031] <= 18'h1e4a1;
	 filter_in_data_log_force[2032] <= 18'h200bb;
	 filter_in_data_log_force[2033] <= 18'h1f3d3;
	 filter_in_data_log_force[2034] <= 18'h23ba6;
	 filter_in_data_log_force[2035] <= 18'h17567;
	 filter_in_data_log_force[2036] <= 18'h2f27e;
	 filter_in_data_log_force[2037] <= 18'h0948e;
	 filter_in_data_log_force[2038] <= 18'h3ecd6;
	 filter_in_data_log_force[2039] <= 18'h39204;
	 filter_in_data_log_force[2040] <= 18'h0e6b4;
	 filter_in_data_log_force[2041] <= 18'h2b030;
	 filter_in_data_log_force[2042] <= 18'h1a381;
	 filter_in_data_log_force[2043] <= 18'h22266;
	 filter_in_data_log_force[2044] <= 18'h1fbb2;
	 filter_in_data_log_force[2045] <= 18'h202e2;
	 filter_in_data_log_force[2046] <= 18'h1e2dc;
	 filter_in_data_log_force[2047] <= 18'h250a2;
	 filter_in_data_log_force[2048] <= 18'h16649;
	 filter_in_data_log_force[2049] <= 18'h2f3d8;
	 filter_in_data_log_force[2050] <= 18'h0a61b;
	 filter_in_data_log_force[2051] <= 18'h3c67b;
	 filter_in_data_log_force[2052] <= 18'h3cbc0;
	 filter_in_data_log_force[2053] <= 18'h09e28;
	 filter_in_data_log_force[2054] <= 18'h30057;
	 filter_in_data_log_force[2055] <= 18'h154e9;
	 filter_in_data_log_force[2056] <= 18'h26525;
	 filter_in_data_log_force[2057] <= 18'h1cf50;
	 filter_in_data_log_force[2058] <= 18'h20f07;
	 filter_in_data_log_force[2059] <= 18'h1ff62;
	 filter_in_data_log_force[2060] <= 18'h20520;
	 filter_in_data_log_force[2061] <= 18'h1e47c;
	 filter_in_data_log_force[2062] <= 18'h2422c;
	 filter_in_data_log_force[2063] <= 18'h188ff;
	 filter_in_data_log_force[2064] <= 18'h2b799;
	 filter_in_data_log_force[2065] <= 18'h0feb1;
	 filter_in_data_log_force[2066] <= 18'h3516a;
	 filter_in_data_log_force[2067] <= 18'h05acf;
	 filter_in_data_log_force[2068] <= 18'h3fa0a;
	 filter_in_data_log_force[2069] <= 18'h3b278;
	 filter_in_data_log_force[2070] <= 18'h09d7c;
	 filter_in_data_log_force[2071] <= 18'h317fe;
	 filter_in_data_log_force[2072] <= 18'h12b88;
	 filter_in_data_log_force[2073] <= 18'h29930;
	 filter_in_data_log_force[2074] <= 18'h198ef;
	 filter_in_data_log_force[2075] <= 18'h23eb2;
	 filter_in_data_log_force[2076] <= 18'h1dfa1;
	 filter_in_data_log_force[2077] <= 18'h20c1c;
	 filter_in_data_log_force[2078] <= 18'h1fe4f;
	 filter_in_data_log_force[2079] <= 18'h200b3;
	 filter_in_data_log_force[2080] <= 18'h1f779;
	 filter_in_data_log_force[2081] <= 18'h21873;
	 filter_in_data_log_force[2082] <= 18'h1d05b;
	 filter_in_data_log_force[2083] <= 18'h24d36;
	 filter_in_data_log_force[2084] <= 18'h18fc6;
	 filter_in_data_log_force[2085] <= 18'h297c1;
	 filter_in_data_log_force[2086] <= 18'h13d21;
	 filter_in_data_log_force[2087] <= 18'h2f0b1;
	 filter_in_data_log_force[2088] <= 18'h0dfa1;
	 filter_in_data_log_force[2089] <= 18'h35122;
	 filter_in_data_log_force[2090] <= 18'h07dbb;
	 filter_in_data_log_force[2091] <= 18'h3b327;
	 filter_in_data_log_force[2092] <= 18'h01cc6;
	 filter_in_data_log_force[2093] <= 18'h01204;
	 filter_in_data_log_force[2094] <= 18'h3c0e0;
	 filter_in_data_log_force[2095] <= 18'h06a3c;
	 filter_in_data_log_force[2096] <= 18'h36ce7;
	 filter_in_data_log_force[2097] <= 18'h0b986;
	 filter_in_data_log_force[2098] <= 18'h3229b;
	 filter_in_data_log_force[2099] <= 18'h0fea3;
	 filter_in_data_log_force[2100] <= 18'h2e2c4;
	 filter_in_data_log_force[2101] <= 18'h13933;
	 filter_in_data_log_force[2102] <= 18'h2ad69;
	 filter_in_data_log_force[2103] <= 18'h00000;
	 filter_in_data_log_force[2104] <= 18'h00000;
	 filter_in_data_log_force[2105] <= 18'h00000;
	 filter_in_data_log_force[2106] <= 18'h00000;
	 filter_in_data_log_force[2107] <= 18'h00000;
	 filter_in_data_log_force[2108] <= 18'h00000;
	 filter_in_data_log_force[2109] <= 18'h00000;
	 filter_in_data_log_force[2110] <= 18'h00000;
	 filter_in_data_log_force[2111] <= 18'h00000;
	 filter_in_data_log_force[2112] <= 18'h00000;
	 filter_in_data_log_force[2113] <= 18'h00000;
	 filter_in_data_log_force[2114] <= 18'h2b8f4;
	 filter_in_data_log_force[2115] <= 18'h22e22;
	 filter_in_data_log_force[2116] <= 18'h0e488;
	 filter_in_data_log_force[2117] <= 18'h363c7;
	 filter_in_data_log_force[2118] <= 18'h0a479;
	 filter_in_data_log_force[2119] <= 18'h38915;
	 filter_in_data_log_force[2120] <= 18'h08267;
	 filter_in_data_log_force[2121] <= 18'h2162b;
	 filter_in_data_log_force[2122] <= 18'h1a46c;
	 filter_in_data_log_force[2123] <= 18'h133c6;
	 filter_in_data_log_force[2124] <= 18'h0fbbf;
	 filter_in_data_log_force[2125] <= 18'h140a1;
	 filter_in_data_log_force[2126] <= 18'h38881;
	 filter_in_data_log_force[2127] <= 18'h07818;
	 filter_in_data_log_force[2128] <= 18'h04d4f;
	 filter_in_data_log_force[2129] <= 18'h01ec6;
	 filter_in_data_log_force[2130] <= 18'h319ac;
	 filter_in_data_log_force[2131] <= 18'h2fe99;
	 filter_in_data_log_force[2132] <= 18'h3ce7a;
	 filter_in_data_log_force[2133] <= 18'h2e92e;
	 filter_in_data_log_force[2134] <= 18'h137c2;
	 filter_in_data_log_force[2135] <= 18'h1f1c5;
	 filter_in_data_log_force[2136] <= 18'h21eb6;
	 filter_in_data_log_force[2137] <= 18'h02485;
	 filter_in_data_log_force[2138] <= 18'h2592b;
	 filter_in_data_log_force[2139] <= 18'h13557;
	 filter_in_data_log_force[2140] <= 18'h1f4e2;
	 filter_in_data_log_force[2141] <= 18'h2448e;
	 filter_in_data_log_force[2142] <= 18'h1c1f2;
	 filter_in_data_log_force[2143] <= 18'h2129d;
	 filter_in_data_log_force[2144] <= 18'h0bc40;
	 filter_in_data_log_force[2145] <= 18'h1228c;
	 filter_in_data_log_force[2146] <= 18'h022f5;
	 filter_in_data_log_force[2147] <= 18'h18a9c;
	 filter_in_data_log_force[2148] <= 18'h19895;
	 filter_in_data_log_force[2149] <= 18'h080f6;
	 filter_in_data_log_force[2150] <= 18'h28d2e;
	 filter_in_data_log_force[2151] <= 18'h2df07;
	 filter_in_data_log_force[2152] <= 18'h2ba83;
	 filter_in_data_log_force[2153] <= 18'h22ad3;
	 filter_in_data_log_force[2154] <= 18'h26d82;
	 filter_in_data_log_force[2155] <= 18'h0773d;
	 filter_in_data_log_force[2156] <= 18'h1c236;
	 filter_in_data_log_force[2157] <= 18'h36af6;
	 filter_in_data_log_force[2158] <= 18'h3a47c;
	 filter_in_data_log_force[2159] <= 18'h1eff9;
	 filter_in_data_log_force[2160] <= 18'h1c846;
	 filter_in_data_log_force[2161] <= 18'h0b4e2;
	 filter_in_data_log_force[2162] <= 18'h1f406;
	 filter_in_data_log_force[2163] <= 18'h1113c;
	 filter_in_data_log_force[2164] <= 18'h358c8;
	 filter_in_data_log_force[2165] <= 18'h0a647;
	 filter_in_data_log_force[2166] <= 18'h2fa06;
	 filter_in_data_log_force[2167] <= 18'h32e99;
	 filter_in_data_log_force[2168] <= 18'h0b881;
	 filter_in_data_log_force[2169] <= 18'h01c84;
	 filter_in_data_log_force[2170] <= 18'h3a579;
	 filter_in_data_log_force[2171] <= 18'h0691a;
	 filter_in_data_log_force[2172] <= 18'h10088;
	 filter_in_data_log_force[2173] <= 18'h0558a;
	 filter_in_data_log_force[2174] <= 18'h03509;
	 filter_in_data_log_force[2175] <= 18'h05594;
	 filter_in_data_log_force[2176] <= 18'h00c1b;
	 filter_in_data_log_force[2177] <= 18'h25493;
	 filter_in_data_log_force[2178] <= 18'h0e0d7;
	 filter_in_data_log_force[2179] <= 18'h1fc10;
	 filter_in_data_log_force[2180] <= 18'h36b0b;
	 filter_in_data_log_force[2181] <= 18'h1e292;
	 filter_in_data_log_force[2182] <= 18'h362c3;
	 filter_in_data_log_force[2183] <= 18'h18bd2;
	 filter_in_data_log_force[2184] <= 18'h3d19c;
	 filter_in_data_log_force[2185] <= 18'h3a759;
	 filter_in_data_log_force[2186] <= 18'h2def5;
	 filter_in_data_log_force[2187] <= 18'h280ac;
	 filter_in_data_log_force[2188] <= 18'h33c54;
	 filter_in_data_log_force[2189] <= 18'h0e788;
	 filter_in_data_log_force[2190] <= 18'h121a9;
	 filter_in_data_log_force[2191] <= 18'h0c670;
	 filter_in_data_log_force[2192] <= 18'h20a0a;
	 filter_in_data_log_force[2193] <= 18'h15f73;
	 filter_in_data_log_force[2194] <= 18'h1b078;
	 filter_in_data_log_force[2195] <= 18'h11575;
	 filter_in_data_log_force[2196] <= 18'h22baf;
	 filter_in_data_log_force[2197] <= 18'h38343;
	 filter_in_data_log_force[2198] <= 18'h0d13e;
	 filter_in_data_log_force[2199] <= 18'h0eb05;
	 filter_in_data_log_force[2200] <= 18'h2e5a9;
	 filter_in_data_log_force[2201] <= 18'h31383;
	 filter_in_data_log_force[2202] <= 18'h0b12f;
	 filter_in_data_log_force[2203] <= 18'h3e8f4;
	 filter_in_data_log_force[2204] <= 18'h07eb0;
	 filter_in_data_log_force[2205] <= 18'h2f21f;
	 filter_in_data_log_force[2206] <= 18'h2b560;
	 filter_in_data_log_force[2207] <= 18'h1518e;
	 filter_in_data_log_force[2208] <= 18'h11154;
	 filter_in_data_log_force[2209] <= 18'h1bce8;
	 filter_in_data_log_force[2210] <= 18'h26e7a;
	 filter_in_data_log_force[2211] <= 18'h2ba9a;
	 filter_in_data_log_force[2212] <= 18'h26579;
	 filter_in_data_log_force[2213] <= 18'h3f585;
	 filter_in_data_log_force[2214] <= 18'h2c5e2;
	 filter_in_data_log_force[2215] <= 18'h19565;
	 filter_in_data_log_force[2216] <= 18'h26578;
	 filter_in_data_log_force[2217] <= 18'h22d3a;
	 filter_in_data_log_force[2218] <= 18'h03aac;
	 filter_in_data_log_force[2219] <= 18'h11709;
	 filter_in_data_log_force[2220] <= 18'h33f6d;
	 filter_in_data_log_force[2221] <= 18'h2b747;
	 filter_in_data_log_force[2222] <= 18'h35b17;
	 filter_in_data_log_force[2223] <= 18'h2d730;
	 filter_in_data_log_force[2224] <= 18'h00a65;
	 filter_in_data_log_force[2225] <= 18'h1a01e;
	 filter_in_data_log_force[2226] <= 18'h08405;
	 filter_in_data_log_force[2227] <= 18'h267f8;
	 filter_in_data_log_force[2228] <= 18'h3903c;
	 filter_in_data_log_force[2229] <= 18'h237ed;
	 filter_in_data_log_force[2230] <= 18'h00150;
	 filter_in_data_log_force[2231] <= 18'h3ba15;
	 filter_in_data_log_force[2232] <= 18'h1fd80;
	 filter_in_data_log_force[2233] <= 18'h13f15;
	 filter_in_data_log_force[2234] <= 18'h3f14f;
	 filter_in_data_log_force[2235] <= 18'h193ea;
	 filter_in_data_log_force[2236] <= 18'h28cd9;
	 filter_in_data_log_force[2237] <= 18'h38f5d;
	 filter_in_data_log_force[2238] <= 18'h1b59d;
	 filter_in_data_log_force[2239] <= 18'h1ab84;
	 filter_in_data_log_force[2240] <= 18'h0dab3;
	 filter_in_data_log_force[2241] <= 18'h0792d;
	 filter_in_data_log_force[2242] <= 18'h35f87;
	 filter_in_data_log_force[2243] <= 18'h1be7e;
	 filter_in_data_log_force[2244] <= 18'h27fc5;
	 filter_in_data_log_force[2245] <= 18'h0ec1f;
	 filter_in_data_log_force[2246] <= 18'h095fe;
	 filter_in_data_log_force[2247] <= 18'h15526;
	 filter_in_data_log_force[2248] <= 18'h397d7;
	 filter_in_data_log_force[2249] <= 18'h0ffd1;
	 filter_in_data_log_force[2250] <= 18'h15744;
	 filter_in_data_log_force[2251] <= 18'h34a33;
	 filter_in_data_log_force[2252] <= 18'h03584;
	 filter_in_data_log_force[2253] <= 18'h1eaa1;
	 filter_in_data_log_force[2254] <= 18'h0327e;
	 filter_in_data_log_force[2255] <= 18'h3525b;
	 filter_in_data_log_force[2256] <= 18'h07a57;
	 filter_in_data_log_force[2257] <= 18'h3714b;
	 filter_in_data_log_force[2258] <= 18'h106aa;
	 filter_in_data_log_force[2259] <= 18'h3a7d6;
	 filter_in_data_log_force[2260] <= 18'h3f829;
	 filter_in_data_log_force[2261] <= 18'h0c76b;
	 filter_in_data_log_force[2262] <= 18'h1e414;
	 filter_in_data_log_force[2263] <= 18'h34f9f;
	 filter_in_data_log_force[2264] <= 18'h159e9;
	 filter_in_data_log_force[2265] <= 18'h0f4cf;
	 filter_in_data_log_force[2266] <= 18'h1d113;
	 filter_in_data_log_force[2267] <= 18'h220b0;
	 filter_in_data_log_force[2268] <= 18'h36d6f;
	 filter_in_data_log_force[2269] <= 18'h0a68f;
	 filter_in_data_log_force[2270] <= 18'h32042;
	 filter_in_data_log_force[2271] <= 18'h2ebea;
	 filter_in_data_log_force[2272] <= 18'h0d832;
	 filter_in_data_log_force[2273] <= 18'h07f90;
	 filter_in_data_log_force[2274] <= 18'h05cc9;
	 filter_in_data_log_force[2275] <= 18'h0a44a;
	 filter_in_data_log_force[2276] <= 18'h230b2;
	 filter_in_data_log_force[2277] <= 18'h36528;
	 filter_in_data_log_force[2278] <= 18'h3ce2c;
	 filter_in_data_log_force[2279] <= 18'h2f6b0;
	 filter_in_data_log_force[2280] <= 18'h0dc35;
	 filter_in_data_log_force[2281] <= 18'h16cbb;
	 filter_in_data_log_force[2282] <= 18'h32044;
	 filter_in_data_log_force[2283] <= 18'h0ec99;
	 filter_in_data_log_force[2284] <= 18'h28d12;
	 filter_in_data_log_force[2285] <= 18'h158ce;
	 filter_in_data_log_force[2286] <= 18'h28dee;
	 filter_in_data_log_force[2287] <= 18'h05a54;
	 filter_in_data_log_force[2288] <= 18'h376f2;
	 filter_in_data_log_force[2289] <= 18'h13a1f;
	 filter_in_data_log_force[2290] <= 18'h003df;
	 filter_in_data_log_force[2291] <= 18'h3f558;
	 filter_in_data_log_force[2292] <= 18'h18219;
	 filter_in_data_log_force[2293] <= 18'h3699e;
	 filter_in_data_log_force[2294] <= 18'h3cc3b;
	 filter_in_data_log_force[2295] <= 18'h1daa8;
	 filter_in_data_log_force[2296] <= 18'h22b50;
	 filter_in_data_log_force[2297] <= 18'h1e44f;
	 filter_in_data_log_force[2298] <= 18'h2c1bf;
	 filter_in_data_log_force[2299] <= 18'h0ab22;
	 filter_in_data_log_force[2300] <= 18'h05884;
	 filter_in_data_log_force[2301] <= 18'h0b351;
	 filter_in_data_log_force[2302] <= 18'h371b0;
	 filter_in_data_log_force[2303] <= 18'h07b2a;
	 filter_in_data_log_force[2304] <= 18'h13e9e;
	 filter_in_data_log_force[2305] <= 18'h213b8;
	 filter_in_data_log_force[2306] <= 18'h255e3;
	 filter_in_data_log_force[2307] <= 18'h1e632;
	 filter_in_data_log_force[2308] <= 18'h09afb;
	 filter_in_data_log_force[2309] <= 18'h2ecca;
	 filter_in_data_log_force[2310] <= 18'h39d2d;
	 filter_in_data_log_force[2311] <= 18'h27cf3;
	 filter_in_data_log_force[2312] <= 18'h312e2;
	 filter_in_data_log_force[2313] <= 18'h30809;
	 filter_in_data_log_force[2314] <= 18'h353a0;
	 filter_in_data_log_force[2315] <= 18'h29be3;
	 filter_in_data_log_force[2316] <= 18'h3645c;
	 filter_in_data_log_force[2317] <= 18'h27c94;
	 filter_in_data_log_force[2318] <= 18'h1895f;
	 filter_in_data_log_force[2319] <= 18'h2608b;
	 filter_in_data_log_force[2320] <= 18'h1b85d;
	 filter_in_data_log_force[2321] <= 18'h39899;
	 filter_in_data_log_force[2322] <= 18'h2308a;
	 filter_in_data_log_force[2323] <= 18'h35e97;
	 filter_in_data_log_force[2324] <= 18'h0f1a1;
	 filter_in_data_log_force[2325] <= 18'h12dc1;
	 filter_in_data_log_force[2326] <= 18'h02dfc;
	 filter_in_data_log_force[2327] <= 18'h0beb1;
	 filter_in_data_log_force[2328] <= 18'h19314;
	 filter_in_data_log_force[2329] <= 18'h2381b;
	 filter_in_data_log_force[2330] <= 18'h336f3;
	 filter_in_data_log_force[2331] <= 18'h22f4d;
	 filter_in_data_log_force[2332] <= 18'h2c82b;
	 filter_in_data_log_force[2333] <= 18'h0e173;
	 filter_in_data_log_force[2334] <= 18'h0e313;
	 filter_in_data_log_force[2335] <= 18'h182de;
	 filter_in_data_log_force[2336] <= 18'h05469;
	 filter_in_data_log_force[2337] <= 18'h24861;
	 filter_in_data_log_force[2338] <= 18'h1b0e4;
	 filter_in_data_log_force[2339] <= 18'h13395;
	 filter_in_data_log_force[2340] <= 18'h324cf;
	 filter_in_data_log_force[2341] <= 18'h02cb6;
	 filter_in_data_log_force[2342] <= 18'h1f069;
	 filter_in_data_log_force[2343] <= 18'h0dcdb;
	 filter_in_data_log_force[2344] <= 18'h15b1b;
	 filter_in_data_log_force[2345] <= 18'h3bba9;
	 filter_in_data_log_force[2346] <= 18'h3e1eb;
	 filter_in_data_log_force[2347] <= 18'h03e2c;
	 filter_in_data_log_force[2348] <= 18'h3138d;
	 filter_in_data_log_force[2349] <= 18'h0feff;
	 filter_in_data_log_force[2350] <= 18'h003fb;
	 filter_in_data_log_force[2351] <= 18'h09655;
	 filter_in_data_log_force[2352] <= 18'h33b22;
	 filter_in_data_log_force[2353] <= 18'h28e0e;
	 filter_in_data_log_force[2354] <= 18'h3e6fd;
	 filter_in_data_log_force[2355] <= 18'h37329;
	 filter_in_data_log_force[2356] <= 18'h12707;
	 filter_in_data_log_force[2357] <= 18'h11f06;
	 filter_in_data_log_force[2358] <= 18'h0ac8e;
	 filter_in_data_log_force[2359] <= 18'h288b5;
	 filter_in_data_log_force[2360] <= 18'h21613;
	 filter_in_data_log_force[2361] <= 18'h03d47;
	 filter_in_data_log_force[2362] <= 18'h3340a;
	 filter_in_data_log_force[2363] <= 18'h1c1f5;
	 filter_in_data_log_force[2364] <= 18'h1ec72;
	 filter_in_data_log_force[2365] <= 18'h32580;
	 filter_in_data_log_force[2366] <= 18'h1340a;
	 filter_in_data_log_force[2367] <= 18'h1959e;
	 filter_in_data_log_force[2368] <= 18'h063de;
	 filter_in_data_log_force[2369] <= 18'h1893c;
	 filter_in_data_log_force[2370] <= 18'h1c662;
	 filter_in_data_log_force[2371] <= 18'h03256;
	 filter_in_data_log_force[2372] <= 18'h0e9de;
	 filter_in_data_log_force[2373] <= 18'h04e9a;
	 filter_in_data_log_force[2374] <= 18'h21a7a;
	 filter_in_data_log_force[2375] <= 18'h3c93f;
	 filter_in_data_log_force[2376] <= 18'h095d0;
	 filter_in_data_log_force[2377] <= 18'h015b6;
	 filter_in_data_log_force[2378] <= 18'h37d40;
	 filter_in_data_log_force[2379] <= 18'h1bfa0;
	 filter_in_data_log_force[2380] <= 18'h15171;
	 filter_in_data_log_force[2381] <= 18'h16577;
	 filter_in_data_log_force[2382] <= 18'h37d7a;
	 filter_in_data_log_force[2383] <= 18'h05f6c;
	 filter_in_data_log_force[2384] <= 18'h17d7e;
	 filter_in_data_log_force[2385] <= 18'h1bbe8;
	 filter_in_data_log_force[2386] <= 18'h0ac82;
	 filter_in_data_log_force[2387] <= 18'h2d3bd;
	 filter_in_data_log_force[2388] <= 18'h09d8b;
	 filter_in_data_log_force[2389] <= 18'h249c8;
	 filter_in_data_log_force[2390] <= 18'h3a07d;
	 filter_in_data_log_force[2391] <= 18'h0aaf0;
	 filter_in_data_log_force[2392] <= 18'h1bc23;
	 filter_in_data_log_force[2393] <= 18'h13e6a;
	 filter_in_data_log_force[2394] <= 18'h3f02d;
	 filter_in_data_log_force[2395] <= 18'h106e9;
	 filter_in_data_log_force[2396] <= 18'h3ab0e;
	 filter_in_data_log_force[2397] <= 18'h1e31c;
	 filter_in_data_log_force[2398] <= 18'h1f3b0;
	 filter_in_data_log_force[2399] <= 18'h174e3;
	 filter_in_data_log_force[2400] <= 18'h38e38;
	 filter_in_data_log_force[2401] <= 18'h3d1a8;
	 filter_in_data_log_force[2402] <= 18'h2fc9c;
	 filter_in_data_log_force[2403] <= 18'h12340;
	 filter_in_data_log_force[2404] <= 18'h18807;
	 filter_in_data_log_force[2405] <= 18'h1a7a4;
	 filter_in_data_log_force[2406] <= 18'h03baf;
	 filter_in_data_log_force[2407] <= 18'h0653e;
	 filter_in_data_log_force[2408] <= 18'h29873;
	 filter_in_data_log_force[2409] <= 18'h1994e;
	 filter_in_data_log_force[2410] <= 18'h3cd34;
	 filter_in_data_log_force[2411] <= 18'h2d29c;
	 filter_in_data_log_force[2412] <= 18'h1993e;
	 filter_in_data_log_force[2413] <= 18'h10ce3;
	 filter_in_data_log_force[2414] <= 18'h187aa;
	 filter_in_data_log_force[2415] <= 18'h323ca;
	 filter_in_data_log_force[2416] <= 18'h0b162;
	 filter_in_data_log_force[2417] <= 18'h0a839;
	 filter_in_data_log_force[2418] <= 18'h27dc3;
	 filter_in_data_log_force[2419] <= 18'h3a118;
	 filter_in_data_log_force[2420] <= 18'h319e5;
	 filter_in_data_log_force[2421] <= 18'h0dddf;
	 filter_in_data_log_force[2422] <= 18'h32230;
	 filter_in_data_log_force[2423] <= 18'h195b5;
	 filter_in_data_log_force[2424] <= 18'h14e6b;
	 filter_in_data_log_force[2425] <= 18'h38f63;
	 filter_in_data_log_force[2426] <= 18'h3fdda;
	 filter_in_data_log_force[2427] <= 18'h0c77b;
	 filter_in_data_log_force[2428] <= 18'h15665;
	 filter_in_data_log_force[2429] <= 18'h07043;
	 filter_in_data_log_force[2430] <= 18'h04c88;
	 filter_in_data_log_force[2431] <= 18'h34dde;
	 filter_in_data_log_force[2432] <= 18'h3d361;
	 filter_in_data_log_force[2433] <= 18'h0daed;
	 filter_in_data_log_force[2434] <= 18'h189a1;
	 filter_in_data_log_force[2435] <= 18'h0e228;
	 filter_in_data_log_force[2436] <= 18'h2130f;
	 filter_in_data_log_force[2437] <= 18'h0b2f9;
	 filter_in_data_log_force[2438] <= 18'h3c108;
	 filter_in_data_log_force[2439] <= 18'h3c054;
	 filter_in_data_log_force[2440] <= 18'h277d9;
	 filter_in_data_log_force[2441] <= 18'h1423c;
	 filter_in_data_log_force[2442] <= 18'h34ca7;
	 filter_in_data_log_force[2443] <= 18'h2fc23;
	 filter_in_data_log_force[2444] <= 18'h35ef0;
	 filter_in_data_log_force[2445] <= 18'h380b5;
	 filter_in_data_log_force[2446] <= 18'h02fac;
	 filter_in_data_log_force[2447] <= 18'h03f68;
	 filter_in_data_log_force[2448] <= 18'h39552;
	 filter_in_data_log_force[2449] <= 18'h397b0;
	 filter_in_data_log_force[2450] <= 18'h00fbc;
	 filter_in_data_log_force[2451] <= 18'h0a150;
	 filter_in_data_log_force[2452] <= 18'h1cdbd;
	 filter_in_data_log_force[2453] <= 18'h0e3af;
	 filter_in_data_log_force[2454] <= 18'h399af;
	 filter_in_data_log_force[2455] <= 18'h153d6;
	 filter_in_data_log_force[2456] <= 18'h28990;
	 filter_in_data_log_force[2457] <= 18'h23deb;
	 filter_in_data_log_force[2458] <= 18'h25645;
	 filter_in_data_log_force[2459] <= 18'h2a7d5;
	 filter_in_data_log_force[2460] <= 18'h34c00;
	 filter_in_data_log_force[2461] <= 18'h334f8;
	 filter_in_data_log_force[2462] <= 18'h20bf6;
	 filter_in_data_log_force[2463] <= 18'h028dd;
	 filter_in_data_log_force[2464] <= 18'h261a9;
	 filter_in_data_log_force[2465] <= 18'h29608;
	 filter_in_data_log_force[2466] <= 18'h0864a;
	 filter_in_data_log_force[2467] <= 18'h16ff2;
	 filter_in_data_log_force[2468] <= 18'h1e59a;
	 filter_in_data_log_force[2469] <= 18'h0488a;
	 filter_in_data_log_force[2470] <= 18'h1fcc6;
	 filter_in_data_log_force[2471] <= 18'h036d4;
	 filter_in_data_log_force[2472] <= 18'h00fd4;
	 filter_in_data_log_force[2473] <= 18'h3529e;
	 filter_in_data_log_force[2474] <= 18'h3b852;
	 filter_in_data_log_force[2475] <= 18'h3f79c;
	 filter_in_data_log_force[2476] <= 18'h248be;
	 filter_in_data_log_force[2477] <= 18'h18d0c;
	 filter_in_data_log_force[2478] <= 18'h2422f;
	 filter_in_data_log_force[2479] <= 18'h3bea7;
	 filter_in_data_log_force[2480] <= 18'h14e78;
	 filter_in_data_log_force[2481] <= 18'h39401;
	 filter_in_data_log_force[2482] <= 18'h07433;
	 filter_in_data_log_force[2483] <= 18'h1464a;
	 filter_in_data_log_force[2484] <= 18'h18b81;
	 filter_in_data_log_force[2485] <= 18'h1b975;
	 filter_in_data_log_force[2486] <= 18'h2c35d;
	 filter_in_data_log_force[2487] <= 18'h308ca;
	 filter_in_data_log_force[2488] <= 18'h1976a;
	 filter_in_data_log_force[2489] <= 18'h05f9a;
	 filter_in_data_log_force[2490] <= 18'h003ef;
	 filter_in_data_log_force[2491] <= 18'h07384;
	 filter_in_data_log_force[2492] <= 18'h14717;
	 filter_in_data_log_force[2493] <= 18'h020a8;
	 filter_in_data_log_force[2494] <= 18'h2ceed;
	 filter_in_data_log_force[2495] <= 18'h3d0c9;
	 filter_in_data_log_force[2496] <= 18'h3b62e;
	 filter_in_data_log_force[2497] <= 18'h1dd3d;
	 filter_in_data_log_force[2498] <= 18'h07af0;
	 filter_in_data_log_force[2499] <= 18'h0c814;
	 filter_in_data_log_force[2500] <= 18'h0e173;
	 filter_in_data_log_force[2501] <= 18'h36338;
	 filter_in_data_log_force[2502] <= 18'h01166;
	 filter_in_data_log_force[2503] <= 18'h03a0e;
	 filter_in_data_log_force[2504] <= 18'h2a040;
	 filter_in_data_log_force[2505] <= 18'h03f8c;
	 filter_in_data_log_force[2506] <= 18'h0c77b;
	 filter_in_data_log_force[2507] <= 18'h3b4b1;
	 filter_in_data_log_force[2508] <= 18'h15857;
	 filter_in_data_log_force[2509] <= 18'h0ecf1;
	 filter_in_data_log_force[2510] <= 18'h370ac;
	 filter_in_data_log_force[2511] <= 18'h3d11d;
	 filter_in_data_log_force[2512] <= 18'h38baa;
	 filter_in_data_log_force[2513] <= 18'h11a2b;
	 filter_in_data_log_force[2514] <= 18'h0efe5;
	 filter_in_data_log_force[2515] <= 18'h3b89b;
	 filter_in_data_log_force[2516] <= 18'h0c667;
	 filter_in_data_log_force[2517] <= 18'h1c7e6;
	 filter_in_data_log_force[2518] <= 18'h1230e;
	 filter_in_data_log_force[2519] <= 18'h0d281;
	 filter_in_data_log_force[2520] <= 18'h26ff5;
	 filter_in_data_log_force[2521] <= 18'h38f4a;
	 filter_in_data_log_force[2522] <= 18'h05d16;
	 filter_in_data_log_force[2523] <= 18'h3d668;
	 filter_in_data_log_force[2524] <= 18'h2338c;
	 filter_in_data_log_force[2525] <= 18'h2ea2d;
	 filter_in_data_log_force[2526] <= 18'h15636;
	 filter_in_data_log_force[2527] <= 18'h21005;
	 filter_in_data_log_force[2528] <= 18'h17471;
	 filter_in_data_log_force[2529] <= 18'h24ff1;
	 filter_in_data_log_force[2530] <= 18'h0ad1a;
	 filter_in_data_log_force[2531] <= 18'h00037;
	 filter_in_data_log_force[2532] <= 18'h2df3a;
	 filter_in_data_log_force[2533] <= 18'h04956;
	 filter_in_data_log_force[2534] <= 18'h27d1f;
	 filter_in_data_log_force[2535] <= 18'h0af46;
	 filter_in_data_log_force[2536] <= 18'h065fa;
	 filter_in_data_log_force[2537] <= 18'h23952;
	 filter_in_data_log_force[2538] <= 18'h239b2;
	 filter_in_data_log_force[2539] <= 18'h29c29;
	 filter_in_data_log_force[2540] <= 18'h21418;
	 filter_in_data_log_force[2541] <= 18'h3bd9f;
	 filter_in_data_log_force[2542] <= 18'h15432;
	 filter_in_data_log_force[2543] <= 18'h07835;
	 filter_in_data_log_force[2544] <= 18'h0149d;
	 filter_in_data_log_force[2545] <= 18'h1749a;
	 filter_in_data_log_force[2546] <= 18'h2640b;
	 filter_in_data_log_force[2547] <= 18'h1a1d8;
	 filter_in_data_log_force[2548] <= 18'h26e9c;
	 filter_in_data_log_force[2549] <= 18'h01168;
	 filter_in_data_log_force[2550] <= 18'h29297;
	 filter_in_data_log_force[2551] <= 18'h03ccc;
	 filter_in_data_log_force[2552] <= 18'h204b1;
	 filter_in_data_log_force[2553] <= 18'h11115;
	 filter_in_data_log_force[2554] <= 18'h16514;
	 filter_in_data_log_force[2555] <= 18'h1aad3;
	 filter_in_data_log_force[2556] <= 18'h1f2a8;
	 filter_in_data_log_force[2557] <= 18'h00542;
	 filter_in_data_log_force[2558] <= 18'h315f0;
	 filter_in_data_log_force[2559] <= 18'h2672b;
	 filter_in_data_log_force[2560] <= 18'h0080a;
	 filter_in_data_log_force[2561] <= 18'h057aa;
	 filter_in_data_log_force[2562] <= 18'h10d32;
	 filter_in_data_log_force[2563] <= 18'h254f4;
	 filter_in_data_log_force[2564] <= 18'h0a579;
	 filter_in_data_log_force[2565] <= 18'h01163;
	 filter_in_data_log_force[2566] <= 18'h2af27;
	 filter_in_data_log_force[2567] <= 18'h1c115;
	 filter_in_data_log_force[2568] <= 18'h05ca8;
	 filter_in_data_log_force[2569] <= 18'h3c336;
	 filter_in_data_log_force[2570] <= 18'h1c486;
	 filter_in_data_log_force[2571] <= 18'h09fa8;
	 filter_in_data_log_force[2572] <= 18'h3cecb;
	 filter_in_data_log_force[2573] <= 18'h15bda;
	 filter_in_data_log_force[2574] <= 18'h02168;
	 filter_in_data_log_force[2575] <= 18'h0372e;
	 filter_in_data_log_force[2576] <= 18'h0b863;
	 filter_in_data_log_force[2577] <= 18'h37801;
	 filter_in_data_log_force[2578] <= 18'h2f509;
	 filter_in_data_log_force[2579] <= 18'h050d1;
	 filter_in_data_log_force[2580] <= 18'h177b1;
	 filter_in_data_log_force[2581] <= 18'h3a08a;
	 filter_in_data_log_force[2582] <= 18'h27351;
	 filter_in_data_log_force[2583] <= 18'h3c680;
	 filter_in_data_log_force[2584] <= 18'h33364;
	 filter_in_data_log_force[2585] <= 18'h39b05;
	 filter_in_data_log_force[2586] <= 18'h1555d;
	 filter_in_data_log_force[2587] <= 18'h39d51;
	 filter_in_data_log_force[2588] <= 18'h38f8a;
	 filter_in_data_log_force[2589] <= 18'h3711a;
	 filter_in_data_log_force[2590] <= 18'h28f9f;
	 filter_in_data_log_force[2591] <= 18'h30a60;
	 filter_in_data_log_force[2592] <= 18'h258e6;
	 filter_in_data_log_force[2593] <= 18'h3b7b4;
	 filter_in_data_log_force[2594] <= 18'h30775;
	 filter_in_data_log_force[2595] <= 18'h330b2;
	 filter_in_data_log_force[2596] <= 18'h3b30e;
	 filter_in_data_log_force[2597] <= 18'h27a11;
	 filter_in_data_log_force[2598] <= 18'h3faf3;
	 filter_in_data_log_force[2599] <= 18'h0d35c;
	 filter_in_data_log_force[2600] <= 18'h2f96b;
	 filter_in_data_log_force[2601] <= 18'h123e9;
	 filter_in_data_log_force[2602] <= 18'h24bde;
	 filter_in_data_log_force[2603] <= 18'h39356;
	 filter_in_data_log_force[2604] <= 18'h2037a;
	 filter_in_data_log_force[2605] <= 18'h2e1f9;
	 filter_in_data_log_force[2606] <= 18'h20155;
	 filter_in_data_log_force[2607] <= 18'h2c1b8;
	 filter_in_data_log_force[2608] <= 18'h291e7;
	 filter_in_data_log_force[2609] <= 18'h31283;
	 filter_in_data_log_force[2610] <= 18'h2b317;
	 filter_in_data_log_force[2611] <= 18'h28dfa;
	 filter_in_data_log_force[2612] <= 18'h06542;
	 filter_in_data_log_force[2613] <= 18'h19aaf;
	 filter_in_data_log_force[2614] <= 18'h1c1ed;
	 filter_in_data_log_force[2615] <= 18'h2e27e;
	 filter_in_data_log_force[2616] <= 18'h3ee41;
	 filter_in_data_log_force[2617] <= 18'h38109;
	 filter_in_data_log_force[2618] <= 18'h0185a;
	 filter_in_data_log_force[2619] <= 18'h30f3b;
	 filter_in_data_log_force[2620] <= 18'h245ff;
	 filter_in_data_log_force[2621] <= 18'h3becd;
	 filter_in_data_log_force[2622] <= 18'h2b207;
	 filter_in_data_log_force[2623] <= 18'h21abc;
	 filter_in_data_log_force[2624] <= 18'h1d197;
	 filter_in_data_log_force[2625] <= 18'h3b8ee;
	 filter_in_data_log_force[2626] <= 18'h1d8a3;
	 filter_in_data_log_force[2627] <= 18'h10cb6;
	 filter_in_data_log_force[2628] <= 18'h20786;
	 filter_in_data_log_force[2629] <= 18'h0b85c;
	 filter_in_data_log_force[2630] <= 18'h0d2e5;
	 filter_in_data_log_force[2631] <= 18'h0949d;
	 filter_in_data_log_force[2632] <= 18'h03591;
	 filter_in_data_log_force[2633] <= 18'h2df58;
	 filter_in_data_log_force[2634] <= 18'h116e7;
	 filter_in_data_log_force[2635] <= 18'h2e980;
	 filter_in_data_log_force[2636] <= 18'h37bc4;
	 filter_in_data_log_force[2637] <= 18'h19050;
	 filter_in_data_log_force[2638] <= 18'h16cee;
	 filter_in_data_log_force[2639] <= 18'h39c18;
	 filter_in_data_log_force[2640] <= 18'h345a7;
	 filter_in_data_log_force[2641] <= 18'h06f3e;
	 filter_in_data_log_force[2642] <= 18'h1a40a;
	 filter_in_data_log_force[2643] <= 18'h1a2eb;
	 filter_in_data_log_force[2644] <= 18'h05dcb;
	 filter_in_data_log_force[2645] <= 18'h3548e;
	 filter_in_data_log_force[2646] <= 18'h1698a;
	 filter_in_data_log_force[2647] <= 18'h3c504;
	 filter_in_data_log_force[2648] <= 18'h19e0f;
	 filter_in_data_log_force[2649] <= 18'h221fa;
	 filter_in_data_log_force[2650] <= 18'h02134;
	 filter_in_data_log_force[2651] <= 18'h0ddb1;
	 filter_in_data_log_force[2652] <= 18'h2b79b;
	 filter_in_data_log_force[2653] <= 18'h3589c;
	 filter_in_data_log_force[2654] <= 18'h2c038;
	 filter_in_data_log_force[2655] <= 18'h349a7;
	 filter_in_data_log_force[2656] <= 18'h39d8d;
	 filter_in_data_log_force[2657] <= 18'h031bb;
	 filter_in_data_log_force[2658] <= 18'h231e9;
	 filter_in_data_log_force[2659] <= 18'h035ff;
	 filter_in_data_log_force[2660] <= 18'h31968;
	 filter_in_data_log_force[2661] <= 18'h2f74c;
	 filter_in_data_log_force[2662] <= 18'h2f8fb;
	 filter_in_data_log_force[2663] <= 18'h29ddc;
	 filter_in_data_log_force[2664] <= 18'h1d35f;
	 filter_in_data_log_force[2665] <= 18'h1be1e;
	 filter_in_data_log_force[2666] <= 18'h1465d;
	 filter_in_data_log_force[2667] <= 18'h0e9bd;
	 filter_in_data_log_force[2668] <= 18'h2b408;
	 filter_in_data_log_force[2669] <= 18'h37105;
	 filter_in_data_log_force[2670] <= 18'h2c152;
	 filter_in_data_log_force[2671] <= 18'h2013a;
	 filter_in_data_log_force[2672] <= 18'h34403;
	 filter_in_data_log_force[2673] <= 18'h0cc68;
	 filter_in_data_log_force[2674] <= 18'h08043;
	 filter_in_data_log_force[2675] <= 18'h02c18;
	 filter_in_data_log_force[2676] <= 18'h3c193;
	 filter_in_data_log_force[2677] <= 18'h32653;
	 filter_in_data_log_force[2678] <= 18'h001b3;
	 filter_in_data_log_force[2679] <= 18'h10bd3;
	 filter_in_data_log_force[2680] <= 18'h10cb5;
	 filter_in_data_log_force[2681] <= 18'h04de2;
	 filter_in_data_log_force[2682] <= 18'h0fd9b;
	 filter_in_data_log_force[2683] <= 18'h09507;
	 filter_in_data_log_force[2684] <= 18'h27e2d;
	 filter_in_data_log_force[2685] <= 18'h00481;
	 filter_in_data_log_force[2686] <= 18'h36398;
	 filter_in_data_log_force[2687] <= 18'h25e5c;
	 filter_in_data_log_force[2688] <= 18'h29766;
	 filter_in_data_log_force[2689] <= 18'h2caed;
	 filter_in_data_log_force[2690] <= 18'h0b068;
	 filter_in_data_log_force[2691] <= 18'h3b9de;
	 filter_in_data_log_force[2692] <= 18'h0c712;
	 filter_in_data_log_force[2693] <= 18'h306f3;
	 filter_in_data_log_force[2694] <= 18'h209fe;
	 filter_in_data_log_force[2695] <= 18'h0210f;
	 filter_in_data_log_force[2696] <= 18'h31e19;
	 filter_in_data_log_force[2697] <= 18'h1c8f1;
	 filter_in_data_log_force[2698] <= 18'h1a033;
	 filter_in_data_log_force[2699] <= 18'h3921c;
	 filter_in_data_log_force[2700] <= 18'h21974;
	 filter_in_data_log_force[2701] <= 18'h0af8d;
	 filter_in_data_log_force[2702] <= 18'h15943;
	 filter_in_data_log_force[2703] <= 18'h1e2d1;
	 filter_in_data_log_force[2704] <= 18'h23a4d;
	 filter_in_data_log_force[2705] <= 18'h3cd22;
	 filter_in_data_log_force[2706] <= 18'h05473;
	 filter_in_data_log_force[2707] <= 18'h0bf1e;
	 filter_in_data_log_force[2708] <= 18'h0e0b3;
	 filter_in_data_log_force[2709] <= 18'h099a4;
	 filter_in_data_log_force[2710] <= 18'h0e85c;
	 filter_in_data_log_force[2711] <= 18'h37ed2;
	 filter_in_data_log_force[2712] <= 18'h0538a;
	 filter_in_data_log_force[2713] <= 18'h276e8;
	 filter_in_data_log_force[2714] <= 18'h23b0a;
	 filter_in_data_log_force[2715] <= 18'h1eb48;
	 filter_in_data_log_force[2716] <= 18'h323a9;
	 filter_in_data_log_force[2717] <= 18'h06141;
	 filter_in_data_log_force[2718] <= 18'h1d941;
	 filter_in_data_log_force[2719] <= 18'h2be3d;
	 filter_in_data_log_force[2720] <= 18'h2c5ac;
	 filter_in_data_log_force[2721] <= 18'h35dd8;
	 filter_in_data_log_force[2722] <= 18'h1bb4a;
	 filter_in_data_log_force[2723] <= 18'h3900b;
	 filter_in_data_log_force[2724] <= 18'h317c6;
	 filter_in_data_log_force[2725] <= 18'h29b98;
	 filter_in_data_log_force[2726] <= 18'h396a4;
	 filter_in_data_log_force[2727] <= 18'h37fb7;
	 filter_in_data_log_force[2728] <= 18'h28643;
	 filter_in_data_log_force[2729] <= 18'h3bd7b;
	 filter_in_data_log_force[2730] <= 18'h25db6;
	 filter_in_data_log_force[2731] <= 18'h07561;
	 filter_in_data_log_force[2732] <= 18'h20b3e;
	 filter_in_data_log_force[2733] <= 18'h04b05;
	 filter_in_data_log_force[2734] <= 18'h128af;
	 filter_in_data_log_force[2735] <= 18'h2f104;
	 filter_in_data_log_force[2736] <= 18'h3cac6;
	 filter_in_data_log_force[2737] <= 18'h04706;
	 filter_in_data_log_force[2738] <= 18'h23ee0;
	 filter_in_data_log_force[2739] <= 18'h3fc33;
	 filter_in_data_log_force[2740] <= 18'h091bb;
	 filter_in_data_log_force[2741] <= 18'h2e293;
	 filter_in_data_log_force[2742] <= 18'h15925;
	 filter_in_data_log_force[2743] <= 18'h1e262;
	 filter_in_data_log_force[2744] <= 18'h162b0;
	 filter_in_data_log_force[2745] <= 18'h00625;
	 filter_in_data_log_force[2746] <= 18'h31d92;
	 filter_in_data_log_force[2747] <= 18'h0fc89;
	 filter_in_data_log_force[2748] <= 18'h2f29e;
	 filter_in_data_log_force[2749] <= 18'h1d452;
	 filter_in_data_log_force[2750] <= 18'h07b25;
	 filter_in_data_log_force[2751] <= 18'h066ab;
	 filter_in_data_log_force[2752] <= 18'h2b0bf;
	 filter_in_data_log_force[2753] <= 18'h25c84;
	 filter_in_data_log_force[2754] <= 18'h30563;
	 filter_in_data_log_force[2755] <= 18'h16f2d;
	 filter_in_data_log_force[2756] <= 18'h1a4ef;
	 filter_in_data_log_force[2757] <= 18'h0cc6d;
	 filter_in_data_log_force[2758] <= 18'h0e696;
	 filter_in_data_log_force[2759] <= 18'h2eb67;
	 filter_in_data_log_force[2760] <= 18'h04de1;
	 filter_in_data_log_force[2761] <= 18'h13e15;
	 filter_in_data_log_force[2762] <= 18'h39d89;
	 filter_in_data_log_force[2763] <= 18'h1f429;
	 filter_in_data_log_force[2764] <= 18'h25c29;
	 filter_in_data_log_force[2765] <= 18'h348a5;
	 filter_in_data_log_force[2766] <= 18'h00baf;
	 filter_in_data_log_force[2767] <= 18'h23e10;
	 filter_in_data_log_force[2768] <= 18'h0e71b;
	 filter_in_data_log_force[2769] <= 18'h039ea;
	 filter_in_data_log_force[2770] <= 18'h01e11;
	 filter_in_data_log_force[2771] <= 18'h151e7;
	 filter_in_data_log_force[2772] <= 18'h16f5f;
	 filter_in_data_log_force[2773] <= 18'h127f7;
	 filter_in_data_log_force[2774] <= 18'h34576;
	 filter_in_data_log_force[2775] <= 18'h3cf0f;
	 filter_in_data_log_force[2776] <= 18'h10248;
	 filter_in_data_log_force[2777] <= 18'h27080;
	 filter_in_data_log_force[2778] <= 18'h27060;
	 filter_in_data_log_force[2779] <= 18'h3145c;
	 filter_in_data_log_force[2780] <= 18'h0193b;
	 filter_in_data_log_force[2781] <= 18'h1e3ff;
	 filter_in_data_log_force[2782] <= 18'h0d775;
	 filter_in_data_log_force[2783] <= 18'h33f58;
	 filter_in_data_log_force[2784] <= 18'h32a74;
	 filter_in_data_log_force[2785] <= 18'h166c4;
	 filter_in_data_log_force[2786] <= 18'h1a587;
	 filter_in_data_log_force[2787] <= 18'h08e9e;
	 filter_in_data_log_force[2788] <= 18'h30580;
	 filter_in_data_log_force[2789] <= 18'h25acb;
	 filter_in_data_log_force[2790] <= 18'h15a60;
	 filter_in_data_log_force[2791] <= 18'h056c0;
	 filter_in_data_log_force[2792] <= 18'h1cadd;
	 filter_in_data_log_force[2793] <= 18'h23e7e;
	 filter_in_data_log_force[2794] <= 18'h056ac;
	 filter_in_data_log_force[2795] <= 18'h323f3;
	 filter_in_data_log_force[2796] <= 18'h14f99;
	 filter_in_data_log_force[2797] <= 18'h2c392;
	 filter_in_data_log_force[2798] <= 18'h3c527;
	 filter_in_data_log_force[2799] <= 18'h392da;
	 filter_in_data_log_force[2800] <= 18'h14e69;
	 filter_in_data_log_force[2801] <= 18'h0b51e;
	 filter_in_data_log_force[2802] <= 18'h2d496;
	 filter_in_data_log_force[2803] <= 18'h345bd;
	 filter_in_data_log_force[2804] <= 18'h28906;
	 filter_in_data_log_force[2805] <= 18'h0af94;
	 filter_in_data_log_force[2806] <= 18'h048b2;
	 filter_in_data_log_force[2807] <= 18'h2add7;
	 filter_in_data_log_force[2808] <= 18'h29733;
	 filter_in_data_log_force[2809] <= 18'h3e781;
	 filter_in_data_log_force[2810] <= 18'h1a1e6;
	 filter_in_data_log_force[2811] <= 18'h0356d;
	 filter_in_data_log_force[2812] <= 18'h221bb;
	 filter_in_data_log_force[2813] <= 18'h23728;
	 filter_in_data_log_force[2814] <= 18'h13862;
	 filter_in_data_log_force[2815] <= 18'h3ce35;
	 filter_in_data_log_force[2816] <= 18'h387d4;
	 filter_in_data_log_force[2817] <= 18'h12898;
	 filter_in_data_log_force[2818] <= 18'h37508;
	 filter_in_data_log_force[2819] <= 18'h02120;
	 filter_in_data_log_force[2820] <= 18'h0d8bd;
	 filter_in_data_log_force[2821] <= 18'h17c64;
	 filter_in_data_log_force[2822] <= 18'h35094;
	 filter_in_data_log_force[2823] <= 18'h099b9;
	 filter_in_data_log_force[2824] <= 18'h1e63b;
	 filter_in_data_log_force[2825] <= 18'h24dca;
	 filter_in_data_log_force[2826] <= 18'h0591c;
	 filter_in_data_log_force[2827] <= 18'h3a7d2;
	 filter_in_data_log_force[2828] <= 18'h33c8e;
	 filter_in_data_log_force[2829] <= 18'h30e2b;
	 filter_in_data_log_force[2830] <= 18'h108fa;
	 filter_in_data_log_force[2831] <= 18'h1fb1a;
	 filter_in_data_log_force[2832] <= 18'h2bf0d;
	 filter_in_data_log_force[2833] <= 18'h11fe5;
	 filter_in_data_log_force[2834] <= 18'h2c87f;
	 filter_in_data_log_force[2835] <= 18'h1f82d;
	 filter_in_data_log_force[2836] <= 18'h13584;
	 filter_in_data_log_force[2837] <= 18'h3b268;
	 filter_in_data_log_force[2838] <= 18'h0ea5b;
	 filter_in_data_log_force[2839] <= 18'h3fe50;
	 filter_in_data_log_force[2840] <= 18'h13c68;
	 filter_in_data_log_force[2841] <= 18'h36d11;
	 filter_in_data_log_force[2842] <= 18'h24b00;
	 filter_in_data_log_force[2843] <= 18'h05d2d;
	 filter_in_data_log_force[2844] <= 18'h1a408;
	 filter_in_data_log_force[2845] <= 18'h2c66b;
	 filter_in_data_log_force[2846] <= 18'h3babf;
	 filter_in_data_log_force[2847] <= 18'h0ff24;
	 filter_in_data_log_force[2848] <= 18'h22820;
	 filter_in_data_log_force[2849] <= 18'h1c909;
	 filter_in_data_log_force[2850] <= 18'h10e00;
	 filter_in_data_log_force[2851] <= 18'h03c3b;
	 filter_in_data_log_force[2852] <= 18'h2bc41;
	 filter_in_data_log_force[2853] <= 18'h3fde6;
	 filter_in_data_log_force[2854] <= 18'h01246;
	 filter_in_data_log_force[2855] <= 18'h1fa1b;
	 filter_in_data_log_force[2856] <= 18'h16b5e;
	 filter_in_data_log_force[2857] <= 18'h1d980;
	 filter_in_data_log_force[2858] <= 18'h0b73c;
	 filter_in_data_log_force[2859] <= 18'h39d2f;
	 filter_in_data_log_force[2860] <= 18'h1bd6b;
	 filter_in_data_log_force[2861] <= 18'h3eafe;
	 filter_in_data_log_force[2862] <= 18'h2ed5b;
	 filter_in_data_log_force[2863] <= 18'h395cd;
	 filter_in_data_log_force[2864] <= 18'h0d200;
	 filter_in_data_log_force[2865] <= 18'h03bf7;
	 filter_in_data_log_force[2866] <= 18'h106ca;
	 filter_in_data_log_force[2867] <= 18'h1fb5f;
	 filter_in_data_log_force[2868] <= 18'h1d988;
	 filter_in_data_log_force[2869] <= 18'h023e9;
	 filter_in_data_log_force[2870] <= 18'h1db01;
	 filter_in_data_log_force[2871] <= 18'h27667;
	 filter_in_data_log_force[2872] <= 18'h234af;
	 filter_in_data_log_force[2873] <= 18'h337a7;
	 filter_in_data_log_force[2874] <= 18'h0521e;
	 filter_in_data_log_force[2875] <= 18'h01fb5;
	 filter_in_data_log_force[2876] <= 18'h19ad6;
	 filter_in_data_log_force[2877] <= 18'h02986;
	 filter_in_data_log_force[2878] <= 18'h3ba59;
	 filter_in_data_log_force[2879] <= 18'h02bb1;
	 filter_in_data_log_force[2880] <= 18'h0d983;
	 filter_in_data_log_force[2881] <= 18'h21113;
	 filter_in_data_log_force[2882] <= 18'h13425;
	 filter_in_data_log_force[2883] <= 18'h291ee;
	 filter_in_data_log_force[2884] <= 18'h3e9f5;
	 filter_in_data_log_force[2885] <= 18'h30700;
	 filter_in_data_log_force[2886] <= 18'h379f3;
	 filter_in_data_log_force[2887] <= 18'h0a5a6;
	 filter_in_data_log_force[2888] <= 18'h2adae;
	 filter_in_data_log_force[2889] <= 18'h31d7a;
	 filter_in_data_log_force[2890] <= 18'h2cafb;
	 filter_in_data_log_force[2891] <= 18'h2c7c1;
	 filter_in_data_log_force[2892] <= 18'h34eaf;
	 filter_in_data_log_force[2893] <= 18'h18577;
	 filter_in_data_log_force[2894] <= 18'h3e269;
	 filter_in_data_log_force[2895] <= 18'h39daa;
	 filter_in_data_log_force[2896] <= 18'h2b788;
	 filter_in_data_log_force[2897] <= 18'h1e02e;
	 filter_in_data_log_force[2898] <= 18'h3a13c;
	 filter_in_data_log_force[2899] <= 18'h160c1;
	 filter_in_data_log_force[2900] <= 18'h07618;
	 filter_in_data_log_force[2901] <= 18'h381a6;
	 filter_in_data_log_force[2902] <= 18'h1823c;
	 filter_in_data_log_force[2903] <= 18'h123b0;
	 filter_in_data_log_force[2904] <= 18'h3dc1d;
	 filter_in_data_log_force[2905] <= 18'h14183;
	 filter_in_data_log_force[2906] <= 18'h19802;
	 filter_in_data_log_force[2907] <= 18'h3b78a;
	 filter_in_data_log_force[2908] <= 18'h3565a;
	 filter_in_data_log_force[2909] <= 18'h062f7;
	 filter_in_data_log_force[2910] <= 18'h19ba3;
	 filter_in_data_log_force[2911] <= 18'h0ceeb;
	 filter_in_data_log_force[2912] <= 18'h38284;
	 filter_in_data_log_force[2913] <= 18'h0f098;
	 filter_in_data_log_force[2914] <= 18'h1d100;
	 filter_in_data_log_force[2915] <= 18'h02bd7;
	 filter_in_data_log_force[2916] <= 18'h02912;
	 filter_in_data_log_force[2917] <= 18'h33e94;
	 filter_in_data_log_force[2918] <= 18'h248f2;
	 filter_in_data_log_force[2919] <= 18'h2ba59;
	 filter_in_data_log_force[2920] <= 18'h25f38;
	 filter_in_data_log_force[2921] <= 18'h3da9d;
	 filter_in_data_log_force[2922] <= 18'h2098e;
	 filter_in_data_log_force[2923] <= 18'h1a8fd;
	 filter_in_data_log_force[2924] <= 18'h0922b;
	 filter_in_data_log_force[2925] <= 18'h20174;
	 filter_in_data_log_force[2926] <= 18'h21f1d;
	 filter_in_data_log_force[2927] <= 18'h2d579;
	 filter_in_data_log_force[2928] <= 18'h3d1e3;
	 filter_in_data_log_force[2929] <= 18'h28252;
	 filter_in_data_log_force[2930] <= 18'h208db;
	 filter_in_data_log_force[2931] <= 18'h0e888;
	 filter_in_data_log_force[2932] <= 18'h36a9e;
	 filter_in_data_log_force[2933] <= 18'h11f2d;
	 filter_in_data_log_force[2934] <= 18'h3bf23;
	 filter_in_data_log_force[2935] <= 18'h3bf08;
	 filter_in_data_log_force[2936] <= 18'h23265;
	 filter_in_data_log_force[2937] <= 18'h232d3;
	 filter_in_data_log_force[2938] <= 18'h25d49;
	 filter_in_data_log_force[2939] <= 18'h0604b;
	 filter_in_data_log_force[2940] <= 18'h2f6df;
	 filter_in_data_log_force[2941] <= 18'h15d90;
	 filter_in_data_log_force[2942] <= 18'h16dc9;
	 filter_in_data_log_force[2943] <= 18'h1dabd;
	 filter_in_data_log_force[2944] <= 18'h3f4a2;
	 filter_in_data_log_force[2945] <= 18'h2e199;
	 filter_in_data_log_force[2946] <= 18'h2e7a3;
	 filter_in_data_log_force[2947] <= 18'h025ac;
	 filter_in_data_log_force[2948] <= 18'h10c66;
	 filter_in_data_log_force[2949] <= 18'h363e9;
	 filter_in_data_log_force[2950] <= 18'h3d84d;
	 filter_in_data_log_force[2951] <= 18'h08eab;
	 filter_in_data_log_force[2952] <= 18'h1ab5a;
	 filter_in_data_log_force[2953] <= 18'h2a573;
	 filter_in_data_log_force[2954] <= 18'h0dcd0;
	 filter_in_data_log_force[2955] <= 18'h04f9b;
	 filter_in_data_log_force[2956] <= 18'h3bbb3;
	 filter_in_data_log_force[2957] <= 18'h18977;
	 filter_in_data_log_force[2958] <= 18'h3927c;
	 filter_in_data_log_force[2959] <= 18'h2b745;
	 filter_in_data_log_force[2960] <= 18'h08889;
	 filter_in_data_log_force[2961] <= 18'h07efa;
	 filter_in_data_log_force[2962] <= 18'h34fd0;
	 filter_in_data_log_force[2963] <= 18'h1363d;
	 filter_in_data_log_force[2964] <= 18'h1ff77;
	 filter_in_data_log_force[2965] <= 18'h1ec86;
	 filter_in_data_log_force[2966] <= 18'h28216;
	 filter_in_data_log_force[2967] <= 18'h2edd0;
	 filter_in_data_log_force[2968] <= 18'h21833;
	 filter_in_data_log_force[2969] <= 18'h06e03;
	 filter_in_data_log_force[2970] <= 18'h27178;
	 filter_in_data_log_force[2971] <= 18'h3a13d;
	 filter_in_data_log_force[2972] <= 18'h1894b;
	 filter_in_data_log_force[2973] <= 18'h0314a;
	 filter_in_data_log_force[2974] <= 18'h379dc;
	 filter_in_data_log_force[2975] <= 18'h2d559;
	 filter_in_data_log_force[2976] <= 18'h3c387;
	 filter_in_data_log_force[2977] <= 18'h1d325;
	 filter_in_data_log_force[2978] <= 18'h27f01;
	 filter_in_data_log_force[2979] <= 18'h3e210;
	 filter_in_data_log_force[2980] <= 18'h16d76;
	 filter_in_data_log_force[2981] <= 18'h22c6f;
	 filter_in_data_log_force[2982] <= 18'h0c439;
	 filter_in_data_log_force[2983] <= 18'h1ea7b;
	 filter_in_data_log_force[2984] <= 18'h32211;
	 filter_in_data_log_force[2985] <= 18'h288fe;
	 filter_in_data_log_force[2986] <= 18'h0bdba;
	 filter_in_data_log_force[2987] <= 18'h1a348;
	 filter_in_data_log_force[2988] <= 18'h07188;
	 filter_in_data_log_force[2989] <= 18'h19995;
	 filter_in_data_log_force[2990] <= 18'h2c613;
	 filter_in_data_log_force[2991] <= 18'h10488;
	 filter_in_data_log_force[2992] <= 18'h36292;
	 filter_in_data_log_force[2993] <= 18'h3acac;
	 filter_in_data_log_force[2994] <= 18'h29f75;
	 filter_in_data_log_force[2995] <= 18'h146a8;
	 filter_in_data_log_force[2996] <= 18'h07fec;
	 filter_in_data_log_force[2997] <= 18'h0f449;
	 filter_in_data_log_force[2998] <= 18'h1386f;
	 filter_in_data_log_force[2999] <= 18'h244d6;
	 filter_in_data_log_force[3000] <= 18'h1cd9c;
	 filter_in_data_log_force[3001] <= 18'h3fd85;
	 filter_in_data_log_force[3002] <= 18'h10545;
	 filter_in_data_log_force[3003] <= 18'h0f839;
	 filter_in_data_log_force[3004] <= 18'h15314;
	 filter_in_data_log_force[3005] <= 18'h2a042;
	 filter_in_data_log_force[3006] <= 18'h3d449;
	 filter_in_data_log_force[3007] <= 18'h078ef;
	 filter_in_data_log_force[3008] <= 18'h1ba8e;
	 filter_in_data_log_force[3009] <= 18'h15721;
	 filter_in_data_log_force[3010] <= 18'h194ea;
	 filter_in_data_log_force[3011] <= 18'h05480;
	 filter_in_data_log_force[3012] <= 18'h054bc;
	 filter_in_data_log_force[3013] <= 18'h16b72;
	 filter_in_data_log_force[3014] <= 18'h223b4;
	 filter_in_data_log_force[3015] <= 18'h18aac;
	 filter_in_data_log_force[3016] <= 18'h3a184;
	 filter_in_data_log_force[3017] <= 18'h22541;
	 filter_in_data_log_force[3018] <= 18'h0fc0e;
	 filter_in_data_log_force[3019] <= 18'h29e8b;
	 filter_in_data_log_force[3020] <= 18'h2935d;
	 filter_in_data_log_force[3021] <= 18'h06c81;
	 filter_in_data_log_force[3022] <= 18'h30497;
	 filter_in_data_log_force[3023] <= 18'h34bef;
	 filter_in_data_log_force[3024] <= 18'h39b6f;
	 filter_in_data_log_force[3025] <= 18'h3a020;
	 filter_in_data_log_force[3026] <= 18'h38b76;
	 filter_in_data_log_force[3027] <= 18'h07070;
	 filter_in_data_log_force[3028] <= 18'h2aae5;
	 filter_in_data_log_force[3029] <= 18'h2c09b;
	 filter_in_data_log_force[3030] <= 18'h260e6;
	 filter_in_data_log_force[3031] <= 18'h34af1;
	 filter_in_data_log_force[3032] <= 18'h11411;
	 filter_in_data_log_force[3033] <= 18'h2efbd;
	 filter_in_data_log_force[3034] <= 18'h0f622;
	 filter_in_data_log_force[3035] <= 18'h0c572;
	 filter_in_data_log_force[3036] <= 18'h14bdb;
	 filter_in_data_log_force[3037] <= 18'h14fd9;
	 filter_in_data_log_force[3038] <= 18'h32c69;
	 filter_in_data_log_force[3039] <= 18'h33ccb;
	 filter_in_data_log_force[3040] <= 18'h01795;
	 filter_in_data_log_force[3041] <= 18'h34d1b;
	 filter_in_data_log_force[3042] <= 18'h153cf;
	 filter_in_data_log_force[3043] <= 18'h13dbe;
	 filter_in_data_log_force[3044] <= 18'h03a5e;
	 filter_in_data_log_force[3045] <= 18'h30d46;
	 filter_in_data_log_force[3046] <= 18'h0b8e6;
	 filter_in_data_log_force[3047] <= 18'h2ef43;
	 filter_in_data_log_force[3048] <= 18'h3d361;
	 filter_in_data_log_force[3049] <= 18'h389cc;
	 filter_in_data_log_force[3050] <= 18'h02787;
	 filter_in_data_log_force[3051] <= 18'h1f781;
	 filter_in_data_log_force[3052] <= 18'h10558;
	 filter_in_data_log_force[3053] <= 18'h1ebfc;
	 filter_in_data_log_force[3054] <= 18'h2f06b;
	 filter_in_data_log_force[3055] <= 18'h01d3f;
	 filter_in_data_log_force[3056] <= 18'h234ac;
	 filter_in_data_log_force[3057] <= 18'h1070a;
	 filter_in_data_log_force[3058] <= 18'h0686d;
	 filter_in_data_log_force[3059] <= 18'h16dbe;
	 filter_in_data_log_force[3060] <= 18'h1f3ff;
	 filter_in_data_log_force[3061] <= 18'h1b7cb;
	 filter_in_data_log_force[3062] <= 18'h3a358;
	 filter_in_data_log_force[3063] <= 18'h2005a;
	 filter_in_data_log_force[3064] <= 18'h029dc;
	 filter_in_data_log_force[3065] <= 18'h2d4b7;
	 filter_in_data_log_force[3066] <= 18'h2e08c;
	 filter_in_data_log_force[3067] <= 18'h34da0;
	 filter_in_data_log_force[3068] <= 18'h26241;
	 filter_in_data_log_force[3069] <= 18'h0fd79;
	 filter_in_data_log_force[3070] <= 18'h0fe79;
	 filter_in_data_log_force[3071] <= 18'h02c57;
	 filter_in_data_log_force[3072] <= 18'h35a3f;
	 filter_in_data_log_force[3073] <= 18'h1544f;
	 filter_in_data_log_force[3074] <= 18'h035d5;
	 filter_in_data_log_force[3075] <= 18'h1d486;
	 filter_in_data_log_force[3076] <= 18'h19243;
	 filter_in_data_log_force[3077] <= 18'h36d0f;
	 filter_in_data_log_force[3078] <= 18'h02f84;
	 filter_in_data_log_force[3079] <= 18'h36301;
	 filter_in_data_log_force[3080] <= 18'h07dc0;
	 filter_in_data_log_force[3081] <= 18'h12fbe;
	 filter_in_data_log_force[3082] <= 18'h0fbc7;
	 filter_in_data_log_force[3083] <= 18'h2808d;
	 filter_in_data_log_force[3084] <= 18'h14a22;
	 filter_in_data_log_force[3085] <= 18'h219c1;
	 filter_in_data_log_force[3086] <= 18'h3a860;
	 filter_in_data_log_force[3087] <= 18'h0ecf6;
	 filter_in_data_log_force[3088] <= 18'h12021;
	 filter_in_data_log_force[3089] <= 18'h3781a;
	 filter_in_data_log_force[3090] <= 18'h0fabf;
	 filter_in_data_log_force[3091] <= 18'h191ae;
	 filter_in_data_log_force[3092] <= 18'h2f86d;
	 filter_in_data_log_force[3093] <= 18'h284b5;
	 filter_in_data_log_force[3094] <= 18'h2e678;
	 filter_in_data_log_force[3095] <= 18'h3666a;
	 filter_in_data_log_force[3096] <= 18'h325fa;
	 filter_in_data_log_force[3097] <= 18'h1b5bf;
	 filter_in_data_log_force[3098] <= 18'h2348c;
	 filter_in_data_log_force[3099] <= 18'h05ee4;
	 filter_in_data_log_force[3100] <= 18'h2a6cf;
	 filter_in_data_log_force[3101] <= 18'h15a87;
	 filter_in_data_log_force[3102] <= 18'h2ab95;
	 filter_in_data_log_force[3103] <= 18'h00241;
	 filter_in_data_log_force[3104] <= 18'h1ff50;
	 filter_in_data_log_force[3105] <= 18'h36bf0;
	 filter_in_data_log_force[3106] <= 18'h23035;
	 filter_in_data_log_force[3107] <= 18'h2daca;
	 filter_in_data_log_force[3108] <= 18'h39763;
	 filter_in_data_log_force[3109] <= 18'h355ad;
	 filter_in_data_log_force[3110] <= 18'h2eb1d;
	 filter_in_data_log_force[3111] <= 18'h1be96;
	 filter_in_data_log_force[3112] <= 18'h0bb96;
	 filter_in_data_log_force[3113] <= 18'h1d934;
	 filter_in_data_log_force[3114] <= 18'h3c07c;
	 filter_in_data_log_force[3115] <= 18'h1c2e8;
	 filter_in_data_log_force[3116] <= 18'h205f9;
	 filter_in_data_log_force[3117] <= 18'h070f4;
	 filter_in_data_log_force[3118] <= 18'h1344d;
	 filter_in_data_log_force[3119] <= 18'h2ee93;
	 filter_in_data_log_force[3120] <= 18'h1bad9;
	 filter_in_data_log_force[3121] <= 18'h10d95;
	 filter_in_data_log_force[3122] <= 18'h14e49;
	 filter_in_data_log_force[3123] <= 18'h04b3a;
	 filter_in_data_log_force[3124] <= 18'h12b9b;
	 filter_in_data_log_force[3125] <= 18'h350f0;
	 filter_in_data_log_force[3126] <= 18'h2e4d3;
	 filter_in_data_log_force[3127] <= 18'h33fe2;
	 filter_in_data_log_force[3128] <= 18'h0568d;
	 filter_in_data_log_force[3129] <= 18'h151d5;
	 filter_in_data_log_force[3130] <= 18'h3296f;
	 filter_in_data_log_force[3131] <= 18'h39c37;
	 filter_in_data_log_force[3132] <= 18'h172bf;
	 filter_in_data_log_force[3133] <= 18'h0757e;
	 filter_in_data_log_force[3134] <= 18'h1f6fa;
	 filter_in_data_log_force[3135] <= 18'h2d096;
	 filter_in_data_log_force[3136] <= 18'h14f10;
	 filter_in_data_log_force[3137] <= 18'h0b415;
	 filter_in_data_log_force[3138] <= 18'h00000;
	 filter_in_data_log_force[3139] <= 18'h00000;
	 filter_in_data_log_force[3140] <= 18'h00000;
	 filter_in_data_log_force[3141] <= 18'h00000;
	 filter_in_data_log_force[3142] <= 18'h00000;
	 filter_in_data_log_force[3143] <= 18'h00000;
	 filter_in_data_log_force[3144] <= 18'h00000;
	 filter_in_data_log_force[3145] <= 18'h00000;
	 filter_in_data_log_force[3146] <= 18'h00000;
	 filter_in_data_log_force[3147] <= 18'h00000;
	 filter_in_data_log_force[3148] <= 18'h00000;

	 // Output data for filter_out
	 filter_out_expected[   0] <= 18'h3d000;
	 filter_out_expected[   1] <= 18'h38000;
	 filter_out_expected[   2] <= 18'h38000;
	 filter_out_expected[   3] <= 18'h00000;
	 filter_out_expected[   4] <= 18'h0b000;
	 filter_out_expected[   5] <= 18'h10000;
	 filter_out_expected[   6] <= 18'h0b000;
	 filter_out_expected[   7] <= 18'h00000;
	 filter_out_expected[   8] <= 18'h38000;
	 filter_out_expected[   9] <= 18'h38000;
	 filter_out_expected[  10] <= 18'h3d000;
	 filter_out_expected[  11] <= 18'h00000;
	 filter_out_expected[  12] <= 18'h00000;
	 filter_out_expected[  13] <= 18'h00000;
	 filter_out_expected[  14] <= 18'h00000;
	 filter_out_expected[  15] <= 18'h00000;
	 filter_out_expected[  16] <= 18'h00000;
	 filter_out_expected[  17] <= 18'h00000;
	 filter_out_expected[  18] <= 18'h00000;
	 filter_out_expected[  19] <= 18'h00000;
	 filter_out_expected[  20] <= 18'h00000;
	 filter_out_expected[  21] <= 18'h00000;
	 filter_out_expected[  22] <= 18'h00000;
	 filter_out_expected[  23] <= 18'h3d000;
	 filter_out_expected[  24] <= 18'h35000;
	 filter_out_expected[  25] <= 18'h2d001;
	 filter_out_expected[  26] <= 18'h2d001;
	 filter_out_expected[  27] <= 18'h38000;
	 filter_out_expected[  28] <= 18'h08000;
	 filter_out_expected[  29] <= 18'h12fff;
	 filter_out_expected[  30] <= 18'h12fff;
	 filter_out_expected[  31] <= 18'h0b000;
	 filter_out_expected[  32] <= 18'h03000;
	 filter_out_expected[  33] <= 18'h03000;
	 filter_out_expected[  34] <= 18'h0b000;
	 filter_out_expected[  35] <= 18'h12fff;
	 filter_out_expected[  36] <= 18'h12fff;
	 filter_out_expected[  37] <= 18'h08000;
	 filter_out_expected[  38] <= 18'h38000;
	 filter_out_expected[  39] <= 18'h2d001;
	 filter_out_expected[  40] <= 18'h2d001;
	 filter_out_expected[  41] <= 18'h35000;
	 filter_out_expected[  42] <= 18'h3d000;
	 filter_out_expected[  43] <= 18'h00000;
	 filter_out_expected[  44] <= 18'h03000;
	 filter_out_expected[  45] <= 18'h0afe8;
	 filter_out_expected[  46] <= 18'h12f90;
	 filter_out_expected[  47] <= 18'h12ef8;
	 filter_out_expected[  48] <= 18'h07e5f;
	 filter_out_expected[  49] <= 18'h37e1f;
	 filter_out_expected[  50] <= 18'h2ce60;
	 filter_out_expected[  51] <= 18'h2cef8;
	 filter_out_expected[  52] <= 18'h34f90;
	 filter_out_expected[  53] <= 18'h3cfe8;
	 filter_out_expected[  54] <= 18'h00000;
	 filter_out_expected[  55] <= 18'h00000;
	 filter_out_expected[  56] <= 18'h00000;
	 filter_out_expected[  57] <= 18'h00000;
	 filter_out_expected[  58] <= 18'h00000;
	 filter_out_expected[  59] <= 18'h00000;
	 filter_out_expected[  60] <= 18'h00000;
	 filter_out_expected[  61] <= 18'h00000;
	 filter_out_expected[  62] <= 18'h00000;
	 filter_out_expected[  63] <= 18'h00000;
	 filter_out_expected[  64] <= 18'h00000;
	 filter_out_expected[  65] <= 18'h00000;
	 filter_out_expected[  66] <= 18'h00000;
	 filter_out_expected[  67] <= 18'h00000;
	 filter_out_expected[  68] <= 18'h00000;
	 filter_out_expected[  69] <= 18'h00000;
	 filter_out_expected[  70] <= 18'h00000;
	 filter_out_expected[  71] <= 18'h00000;
	 filter_out_expected[  72] <= 18'h00000;
	 filter_out_expected[  73] <= 18'h00000;
	 filter_out_expected[  74] <= 18'h00000;
	 filter_out_expected[  75] <= 18'h00000;
	 filter_out_expected[  76] <= 18'h00000;
	 filter_out_expected[  77] <= 18'h00000;
	 filter_out_expected[  78] <= 18'h00000;
	 filter_out_expected[  79] <= 18'h00000;
	 filter_out_expected[  80] <= 18'h00000;
	 filter_out_expected[  81] <= 18'h00000;
	 filter_out_expected[  82] <= 18'h00000;
	 filter_out_expected[  83] <= 18'h00000;
	 filter_out_expected[  84] <= 18'h00000;
	 filter_out_expected[  85] <= 18'h00000;
	 filter_out_expected[  86] <= 18'h00000;
	 filter_out_expected[  87] <= 18'h00000;
	 filter_out_expected[  88] <= 18'h00000;
	 filter_out_expected[  89] <= 18'h00000;
	 filter_out_expected[  90] <= 18'h00000;
	 filter_out_expected[  91] <= 18'h00000;
	 filter_out_expected[  92] <= 18'h00000;
	 filter_out_expected[  93] <= 18'h00000;
	 filter_out_expected[  94] <= 18'h00000;
	 filter_out_expected[  95] <= 18'h00000;
	 filter_out_expected[  96] <= 18'h00000;
	 filter_out_expected[  97] <= 18'h00000;
	 filter_out_expected[  98] <= 18'h00000;
	 filter_out_expected[  99] <= 18'h00000;
	 filter_out_expected[ 100] <= 18'h00000;
	 filter_out_expected[ 101] <= 18'h00000;
	 filter_out_expected[ 102] <= 18'h00000;
	 filter_out_expected[ 103] <= 18'h00000;
	 filter_out_expected[ 104] <= 18'h00000;
	 filter_out_expected[ 105] <= 18'h00000;
	 filter_out_expected[ 106] <= 18'h00000;
	 filter_out_expected[ 107] <= 18'h00000;
	 filter_out_expected[ 108] <= 18'h00000;
	 filter_out_expected[ 109] <= 18'h00000;
	 filter_out_expected[ 110] <= 18'h00000;
	 filter_out_expected[ 111] <= 18'h00000;
	 filter_out_expected[ 112] <= 18'h00000;
	 filter_out_expected[ 113] <= 18'h00000;
	 filter_out_expected[ 114] <= 18'h00000;
	 filter_out_expected[ 115] <= 18'h00000;
	 filter_out_expected[ 116] <= 18'h00000;
	 filter_out_expected[ 117] <= 18'h00000;
	 filter_out_expected[ 118] <= 18'h00000;
	 filter_out_expected[ 119] <= 18'h00000;
	 filter_out_expected[ 120] <= 18'h00000;
	 filter_out_expected[ 121] <= 18'h00000;
	 filter_out_expected[ 122] <= 18'h00000;
	 filter_out_expected[ 123] <= 18'h00000;
	 filter_out_expected[ 124] <= 18'h00000;
	 filter_out_expected[ 125] <= 18'h00000;
	 filter_out_expected[ 126] <= 18'h00000;
	 filter_out_expected[ 127] <= 18'h00000;
	 filter_out_expected[ 128] <= 18'h00000;
	 filter_out_expected[ 129] <= 18'h00000;
	 filter_out_expected[ 130] <= 18'h00000;
	 filter_out_expected[ 131] <= 18'h00000;
	 filter_out_expected[ 132] <= 18'h00000;
	 filter_out_expected[ 133] <= 18'h00000;
	 filter_out_expected[ 134] <= 18'h00000;
	 filter_out_expected[ 135] <= 18'h00000;
	 filter_out_expected[ 136] <= 18'h00000;
	 filter_out_expected[ 137] <= 18'h00000;
	 filter_out_expected[ 138] <= 18'h00000;
	 filter_out_expected[ 139] <= 18'h00000;
	 filter_out_expected[ 140] <= 18'h00000;
	 filter_out_expected[ 141] <= 18'h00000;
	 filter_out_expected[ 142] <= 18'h00000;
	 filter_out_expected[ 143] <= 18'h00000;
	 filter_out_expected[ 144] <= 18'h00000;
	 filter_out_expected[ 145] <= 18'h00000;
	 filter_out_expected[ 146] <= 18'h00000;
	 filter_out_expected[ 147] <= 18'h00000;
	 filter_out_expected[ 148] <= 18'h00000;
	 filter_out_expected[ 149] <= 18'h00000;
	 filter_out_expected[ 150] <= 18'h00000;
	 filter_out_expected[ 151] <= 18'h00000;
	 filter_out_expected[ 152] <= 18'h00000;
	 filter_out_expected[ 153] <= 18'h00000;
	 filter_out_expected[ 154] <= 18'h00000;
	 filter_out_expected[ 155] <= 18'h00000;
	 filter_out_expected[ 156] <= 18'h00000;
	 filter_out_expected[ 157] <= 18'h00000;
	 filter_out_expected[ 158] <= 18'h00000;
	 filter_out_expected[ 159] <= 18'h00000;
	 filter_out_expected[ 160] <= 18'h00000;
	 filter_out_expected[ 161] <= 18'h00000;
	 filter_out_expected[ 162] <= 18'h00000;
	 filter_out_expected[ 163] <= 18'h00000;
	 filter_out_expected[ 164] <= 18'h00000;
	 filter_out_expected[ 165] <= 18'h00000;
	 filter_out_expected[ 166] <= 18'h00000;
	 filter_out_expected[ 167] <= 18'h00000;
	 filter_out_expected[ 168] <= 18'h00000;
	 filter_out_expected[ 169] <= 18'h00000;
	 filter_out_expected[ 170] <= 18'h00000;
	 filter_out_expected[ 171] <= 18'h00000;
	 filter_out_expected[ 172] <= 18'h00000;
	 filter_out_expected[ 173] <= 18'h00000;
	 filter_out_expected[ 174] <= 18'h00000;
	 filter_out_expected[ 175] <= 18'h00000;
	 filter_out_expected[ 176] <= 18'h00000;
	 filter_out_expected[ 177] <= 18'h00000;
	 filter_out_expected[ 178] <= 18'h00000;
	 filter_out_expected[ 179] <= 18'h00000;
	 filter_out_expected[ 180] <= 18'h00000;
	 filter_out_expected[ 181] <= 18'h00000;
	 filter_out_expected[ 182] <= 18'h00000;
	 filter_out_expected[ 183] <= 18'h00000;
	 filter_out_expected[ 184] <= 18'h00000;
	 filter_out_expected[ 185] <= 18'h00000;
	 filter_out_expected[ 186] <= 18'h00000;
	 filter_out_expected[ 187] <= 18'h00000;
	 filter_out_expected[ 188] <= 18'h00000;
	 filter_out_expected[ 189] <= 18'h00000;
	 filter_out_expected[ 190] <= 18'h00000;
	 filter_out_expected[ 191] <= 18'h00000;
	 filter_out_expected[ 192] <= 18'h00000;
	 filter_out_expected[ 193] <= 18'h00000;
	 filter_out_expected[ 194] <= 18'h00000;
	 filter_out_expected[ 195] <= 18'h00000;
	 filter_out_expected[ 196] <= 18'h00000;
	 filter_out_expected[ 197] <= 18'h00000;
	 filter_out_expected[ 198] <= 18'h00000;
	 filter_out_expected[ 199] <= 18'h00000;
	 filter_out_expected[ 200] <= 18'h00000;
	 filter_out_expected[ 201] <= 18'h00000;
	 filter_out_expected[ 202] <= 18'h00000;
	 filter_out_expected[ 203] <= 18'h00000;
	 filter_out_expected[ 204] <= 18'h00000;
	 filter_out_expected[ 205] <= 18'h00000;
	 filter_out_expected[ 206] <= 18'h00000;
	 filter_out_expected[ 207] <= 18'h00000;
	 filter_out_expected[ 208] <= 18'h00000;
	 filter_out_expected[ 209] <= 18'h00000;
	 filter_out_expected[ 210] <= 18'h00000;
	 filter_out_expected[ 211] <= 18'h00000;
	 filter_out_expected[ 212] <= 18'h00000;
	 filter_out_expected[ 213] <= 18'h00000;
	 filter_out_expected[ 214] <= 18'h00000;
	 filter_out_expected[ 215] <= 18'h00000;
	 filter_out_expected[ 216] <= 18'h00000;
	 filter_out_expected[ 217] <= 18'h00000;
	 filter_out_expected[ 218] <= 18'h00000;
	 filter_out_expected[ 219] <= 18'h00000;
	 filter_out_expected[ 220] <= 18'h00000;
	 filter_out_expected[ 221] <= 18'h00000;
	 filter_out_expected[ 222] <= 18'h00000;
	 filter_out_expected[ 223] <= 18'h00000;
	 filter_out_expected[ 224] <= 18'h00000;
	 filter_out_expected[ 225] <= 18'h00000;
	 filter_out_expected[ 226] <= 18'h00000;
	 filter_out_expected[ 227] <= 18'h00000;
	 filter_out_expected[ 228] <= 18'h00000;
	 filter_out_expected[ 229] <= 18'h00000;
	 filter_out_expected[ 230] <= 18'h00000;
	 filter_out_expected[ 231] <= 18'h00000;
	 filter_out_expected[ 232] <= 18'h00000;
	 filter_out_expected[ 233] <= 18'h00000;
	 filter_out_expected[ 234] <= 18'h00000;
	 filter_out_expected[ 235] <= 18'h00000;
	 filter_out_expected[ 236] <= 18'h00000;
	 filter_out_expected[ 237] <= 18'h00000;
	 filter_out_expected[ 238] <= 18'h00000;
	 filter_out_expected[ 239] <= 18'h00000;
	 filter_out_expected[ 240] <= 18'h00000;
	 filter_out_expected[ 241] <= 18'h00000;
	 filter_out_expected[ 242] <= 18'h00000;
	 filter_out_expected[ 243] <= 18'h00000;
	 filter_out_expected[ 244] <= 18'h00000;
	 filter_out_expected[ 245] <= 18'h00000;
	 filter_out_expected[ 246] <= 18'h00000;
	 filter_out_expected[ 247] <= 18'h00000;
	 filter_out_expected[ 248] <= 18'h00000;
	 filter_out_expected[ 249] <= 18'h00000;
	 filter_out_expected[ 250] <= 18'h00000;
	 filter_out_expected[ 251] <= 18'h00000;
	 filter_out_expected[ 252] <= 18'h00000;
	 filter_out_expected[ 253] <= 18'h00000;
	 filter_out_expected[ 254] <= 18'h00000;
	 filter_out_expected[ 255] <= 18'h00000;
	 filter_out_expected[ 256] <= 18'h00000;
	 filter_out_expected[ 257] <= 18'h00000;
	 filter_out_expected[ 258] <= 18'h00000;
	 filter_out_expected[ 259] <= 18'h00000;
	 filter_out_expected[ 260] <= 18'h00000;
	 filter_out_expected[ 261] <= 18'h00000;
	 filter_out_expected[ 262] <= 18'h00000;
	 filter_out_expected[ 263] <= 18'h00000;
	 filter_out_expected[ 264] <= 18'h00000;
	 filter_out_expected[ 265] <= 18'h00000;
	 filter_out_expected[ 266] <= 18'h00000;
	 filter_out_expected[ 267] <= 18'h00000;
	 filter_out_expected[ 268] <= 18'h00000;
	 filter_out_expected[ 269] <= 18'h00000;
	 filter_out_expected[ 270] <= 18'h00000;
	 filter_out_expected[ 271] <= 18'h00000;
	 filter_out_expected[ 272] <= 18'h00000;
	 filter_out_expected[ 273] <= 18'h00000;
	 filter_out_expected[ 274] <= 18'h00000;
	 filter_out_expected[ 275] <= 18'h00000;
	 filter_out_expected[ 276] <= 18'h00000;
	 filter_out_expected[ 277] <= 18'h00000;
	 filter_out_expected[ 278] <= 18'h00000;
	 filter_out_expected[ 279] <= 18'h00000;
	 filter_out_expected[ 280] <= 18'h00000;
	 filter_out_expected[ 281] <= 18'h00000;
	 filter_out_expected[ 282] <= 18'h00000;
	 filter_out_expected[ 283] <= 18'h00000;
	 filter_out_expected[ 284] <= 18'h00000;
	 filter_out_expected[ 285] <= 18'h00000;
	 filter_out_expected[ 286] <= 18'h00000;
	 filter_out_expected[ 287] <= 18'h00000;
	 filter_out_expected[ 288] <= 18'h00000;
	 filter_out_expected[ 289] <= 18'h00000;
	 filter_out_expected[ 290] <= 18'h00000;
	 filter_out_expected[ 291] <= 18'h00000;
	 filter_out_expected[ 292] <= 18'h00000;
	 filter_out_expected[ 293] <= 18'h00000;
	 filter_out_expected[ 294] <= 18'h00000;
	 filter_out_expected[ 295] <= 18'h00000;
	 filter_out_expected[ 296] <= 18'h00000;
	 filter_out_expected[ 297] <= 18'h00000;
	 filter_out_expected[ 298] <= 18'h00000;
	 filter_out_expected[ 299] <= 18'h00000;
	 filter_out_expected[ 300] <= 18'h00000;
	 filter_out_expected[ 301] <= 18'h00000;
	 filter_out_expected[ 302] <= 18'h00000;
	 filter_out_expected[ 303] <= 18'h00000;
	 filter_out_expected[ 304] <= 18'h00000;
	 filter_out_expected[ 305] <= 18'h00000;
	 filter_out_expected[ 306] <= 18'h00000;
	 filter_out_expected[ 307] <= 18'h00000;
	 filter_out_expected[ 308] <= 18'h00000;
	 filter_out_expected[ 309] <= 18'h00000;
	 filter_out_expected[ 310] <= 18'h00000;
	 filter_out_expected[ 311] <= 18'h00000;
	 filter_out_expected[ 312] <= 18'h00000;
	 filter_out_expected[ 313] <= 18'h00000;
	 filter_out_expected[ 314] <= 18'h00000;
	 filter_out_expected[ 315] <= 18'h00000;
	 filter_out_expected[ 316] <= 18'h00000;
	 filter_out_expected[ 317] <= 18'h00000;
	 filter_out_expected[ 318] <= 18'h00000;
	 filter_out_expected[ 319] <= 18'h00000;
	 filter_out_expected[ 320] <= 18'h00000;
	 filter_out_expected[ 321] <= 18'h00000;
	 filter_out_expected[ 322] <= 18'h00000;
	 filter_out_expected[ 323] <= 18'h00000;
	 filter_out_expected[ 324] <= 18'h00000;
	 filter_out_expected[ 325] <= 18'h00000;
	 filter_out_expected[ 326] <= 18'h00000;
	 filter_out_expected[ 327] <= 18'h00000;
	 filter_out_expected[ 328] <= 18'h00000;
	 filter_out_expected[ 329] <= 18'h00000;
	 filter_out_expected[ 330] <= 18'h00000;
	 filter_out_expected[ 331] <= 18'h00000;
	 filter_out_expected[ 332] <= 18'h00000;
	 filter_out_expected[ 333] <= 18'h00000;
	 filter_out_expected[ 334] <= 18'h00000;
	 filter_out_expected[ 335] <= 18'h00000;
	 filter_out_expected[ 336] <= 18'h00000;
	 filter_out_expected[ 337] <= 18'h00000;
	 filter_out_expected[ 338] <= 18'h00000;
	 filter_out_expected[ 339] <= 18'h00000;
	 filter_out_expected[ 340] <= 18'h00000;
	 filter_out_expected[ 341] <= 18'h00000;
	 filter_out_expected[ 342] <= 18'h00000;
	 filter_out_expected[ 343] <= 18'h00000;
	 filter_out_expected[ 344] <= 18'h00000;
	 filter_out_expected[ 345] <= 18'h00000;
	 filter_out_expected[ 346] <= 18'h00000;
	 filter_out_expected[ 347] <= 18'h00000;
	 filter_out_expected[ 348] <= 18'h00000;
	 filter_out_expected[ 349] <= 18'h00000;
	 filter_out_expected[ 350] <= 18'h00000;
	 filter_out_expected[ 351] <= 18'h00000;
	 filter_out_expected[ 352] <= 18'h00000;
	 filter_out_expected[ 353] <= 18'h00000;
	 filter_out_expected[ 354] <= 18'h00000;
	 filter_out_expected[ 355] <= 18'h00000;
	 filter_out_expected[ 356] <= 18'h00000;
	 filter_out_expected[ 357] <= 18'h00000;
	 filter_out_expected[ 358] <= 18'h00000;
	 filter_out_expected[ 359] <= 18'h00000;
	 filter_out_expected[ 360] <= 18'h00000;
	 filter_out_expected[ 361] <= 18'h00000;
	 filter_out_expected[ 362] <= 18'h00000;
	 filter_out_expected[ 363] <= 18'h00000;
	 filter_out_expected[ 364] <= 18'h00000;
	 filter_out_expected[ 365] <= 18'h00000;
	 filter_out_expected[ 366] <= 18'h00000;
	 filter_out_expected[ 367] <= 18'h00000;
	 filter_out_expected[ 368] <= 18'h00000;
	 filter_out_expected[ 369] <= 18'h00000;
	 filter_out_expected[ 370] <= 18'h00000;
	 filter_out_expected[ 371] <= 18'h00000;
	 filter_out_expected[ 372] <= 18'h00000;
	 filter_out_expected[ 373] <= 18'h00000;
	 filter_out_expected[ 374] <= 18'h00000;
	 filter_out_expected[ 375] <= 18'h00000;
	 filter_out_expected[ 376] <= 18'h00000;
	 filter_out_expected[ 377] <= 18'h00000;
	 filter_out_expected[ 378] <= 18'h00000;
	 filter_out_expected[ 379] <= 18'h00000;
	 filter_out_expected[ 380] <= 18'h00000;
	 filter_out_expected[ 381] <= 18'h00000;
	 filter_out_expected[ 382] <= 18'h00000;
	 filter_out_expected[ 383] <= 18'h00000;
	 filter_out_expected[ 384] <= 18'h00000;
	 filter_out_expected[ 385] <= 18'h00000;
	 filter_out_expected[ 386] <= 18'h00000;
	 filter_out_expected[ 387] <= 18'h00000;
	 filter_out_expected[ 388] <= 18'h00000;
	 filter_out_expected[ 389] <= 18'h00000;
	 filter_out_expected[ 390] <= 18'h00000;
	 filter_out_expected[ 391] <= 18'h00000;
	 filter_out_expected[ 392] <= 18'h00000;
	 filter_out_expected[ 393] <= 18'h00000;
	 filter_out_expected[ 394] <= 18'h00000;
	 filter_out_expected[ 395] <= 18'h00000;
	 filter_out_expected[ 396] <= 18'h00000;
	 filter_out_expected[ 397] <= 18'h00000;
	 filter_out_expected[ 398] <= 18'h00000;
	 filter_out_expected[ 399] <= 18'h00000;
	 filter_out_expected[ 400] <= 18'h00000;
	 filter_out_expected[ 401] <= 18'h00000;
	 filter_out_expected[ 402] <= 18'h00000;
	 filter_out_expected[ 403] <= 18'h00000;
	 filter_out_expected[ 404] <= 18'h00000;
	 filter_out_expected[ 405] <= 18'h00000;
	 filter_out_expected[ 406] <= 18'h00000;
	 filter_out_expected[ 407] <= 18'h00000;
	 filter_out_expected[ 408] <= 18'h00000;
	 filter_out_expected[ 409] <= 18'h00000;
	 filter_out_expected[ 410] <= 18'h00000;
	 filter_out_expected[ 411] <= 18'h00000;
	 filter_out_expected[ 412] <= 18'h00000;
	 filter_out_expected[ 413] <= 18'h00000;
	 filter_out_expected[ 414] <= 18'h00000;
	 filter_out_expected[ 415] <= 18'h00000;
	 filter_out_expected[ 416] <= 18'h00000;
	 filter_out_expected[ 417] <= 18'h00000;
	 filter_out_expected[ 418] <= 18'h00000;
	 filter_out_expected[ 419] <= 18'h00000;
	 filter_out_expected[ 420] <= 18'h00000;
	 filter_out_expected[ 421] <= 18'h00000;
	 filter_out_expected[ 422] <= 18'h00000;
	 filter_out_expected[ 423] <= 18'h00000;
	 filter_out_expected[ 424] <= 18'h00000;
	 filter_out_expected[ 425] <= 18'h00000;
	 filter_out_expected[ 426] <= 18'h00000;
	 filter_out_expected[ 427] <= 18'h00000;
	 filter_out_expected[ 428] <= 18'h00000;
	 filter_out_expected[ 429] <= 18'h00000;
	 filter_out_expected[ 430] <= 18'h00000;
	 filter_out_expected[ 431] <= 18'h00000;
	 filter_out_expected[ 432] <= 18'h00000;
	 filter_out_expected[ 433] <= 18'h00000;
	 filter_out_expected[ 434] <= 18'h00000;
	 filter_out_expected[ 435] <= 18'h00000;
	 filter_out_expected[ 436] <= 18'h00000;
	 filter_out_expected[ 437] <= 18'h00000;
	 filter_out_expected[ 438] <= 18'h00000;
	 filter_out_expected[ 439] <= 18'h00000;
	 filter_out_expected[ 440] <= 18'h00000;
	 filter_out_expected[ 441] <= 18'h00000;
	 filter_out_expected[ 442] <= 18'h00000;
	 filter_out_expected[ 443] <= 18'h00000;
	 filter_out_expected[ 444] <= 18'h00000;
	 filter_out_expected[ 445] <= 18'h00000;
	 filter_out_expected[ 446] <= 18'h00000;
	 filter_out_expected[ 447] <= 18'h00000;
	 filter_out_expected[ 448] <= 18'h00000;
	 filter_out_expected[ 449] <= 18'h00000;
	 filter_out_expected[ 450] <= 18'h00000;
	 filter_out_expected[ 451] <= 18'h00000;
	 filter_out_expected[ 452] <= 18'h00000;
	 filter_out_expected[ 453] <= 18'h00000;
	 filter_out_expected[ 454] <= 18'h00000;
	 filter_out_expected[ 455] <= 18'h00000;
	 filter_out_expected[ 456] <= 18'h00000;
	 filter_out_expected[ 457] <= 18'h00000;
	 filter_out_expected[ 458] <= 18'h00000;
	 filter_out_expected[ 459] <= 18'h00000;
	 filter_out_expected[ 460] <= 18'h00000;
	 filter_out_expected[ 461] <= 18'h00000;
	 filter_out_expected[ 462] <= 18'h00000;
	 filter_out_expected[ 463] <= 18'h00000;
	 filter_out_expected[ 464] <= 18'h00000;
	 filter_out_expected[ 465] <= 18'h00000;
	 filter_out_expected[ 466] <= 18'h00000;
	 filter_out_expected[ 467] <= 18'h00000;
	 filter_out_expected[ 468] <= 18'h00000;
	 filter_out_expected[ 469] <= 18'h00000;
	 filter_out_expected[ 470] <= 18'h00000;
	 filter_out_expected[ 471] <= 18'h00000;
	 filter_out_expected[ 472] <= 18'h00000;
	 filter_out_expected[ 473] <= 18'h00000;
	 filter_out_expected[ 474] <= 18'h00000;
	 filter_out_expected[ 475] <= 18'h00000;
	 filter_out_expected[ 476] <= 18'h00000;
	 filter_out_expected[ 477] <= 18'h00000;
	 filter_out_expected[ 478] <= 18'h00000;
	 filter_out_expected[ 479] <= 18'h00000;
	 filter_out_expected[ 480] <= 18'h00000;
	 filter_out_expected[ 481] <= 18'h00000;
	 filter_out_expected[ 482] <= 18'h00000;
	 filter_out_expected[ 483] <= 18'h00000;
	 filter_out_expected[ 484] <= 18'h00000;
	 filter_out_expected[ 485] <= 18'h00000;
	 filter_out_expected[ 486] <= 18'h00000;
	 filter_out_expected[ 487] <= 18'h00000;
	 filter_out_expected[ 488] <= 18'h00000;
	 filter_out_expected[ 489] <= 18'h00000;
	 filter_out_expected[ 490] <= 18'h00000;
	 filter_out_expected[ 491] <= 18'h00000;
	 filter_out_expected[ 492] <= 18'h00000;
	 filter_out_expected[ 493] <= 18'h00000;
	 filter_out_expected[ 494] <= 18'h00000;
	 filter_out_expected[ 495] <= 18'h00000;
	 filter_out_expected[ 496] <= 18'h00000;
	 filter_out_expected[ 497] <= 18'h00000;
	 filter_out_expected[ 498] <= 18'h00000;
	 filter_out_expected[ 499] <= 18'h00000;
	 filter_out_expected[ 500] <= 18'h00000;
	 filter_out_expected[ 501] <= 18'h00000;
	 filter_out_expected[ 502] <= 18'h00000;
	 filter_out_expected[ 503] <= 18'h00000;
	 filter_out_expected[ 504] <= 18'h00000;
	 filter_out_expected[ 505] <= 18'h00000;
	 filter_out_expected[ 506] <= 18'h00000;
	 filter_out_expected[ 507] <= 18'h00000;
	 filter_out_expected[ 508] <= 18'h00000;
	 filter_out_expected[ 509] <= 18'h00000;
	 filter_out_expected[ 510] <= 18'h00000;
	 filter_out_expected[ 511] <= 18'h00000;
	 filter_out_expected[ 512] <= 18'h00000;
	 filter_out_expected[ 513] <= 18'h00000;
	 filter_out_expected[ 514] <= 18'h00000;
	 filter_out_expected[ 515] <= 18'h00000;
	 filter_out_expected[ 516] <= 18'h00000;
	 filter_out_expected[ 517] <= 18'h00000;
	 filter_out_expected[ 518] <= 18'h00000;
	 filter_out_expected[ 519] <= 18'h00000;
	 filter_out_expected[ 520] <= 18'h00000;
	 filter_out_expected[ 521] <= 18'h00000;
	 filter_out_expected[ 522] <= 18'h00000;
	 filter_out_expected[ 523] <= 18'h00000;
	 filter_out_expected[ 524] <= 18'h00000;
	 filter_out_expected[ 525] <= 18'h00000;
	 filter_out_expected[ 526] <= 18'h00000;
	 filter_out_expected[ 527] <= 18'h00000;
	 filter_out_expected[ 528] <= 18'h00000;
	 filter_out_expected[ 529] <= 18'h00000;
	 filter_out_expected[ 530] <= 18'h00000;
	 filter_out_expected[ 531] <= 18'h00000;
	 filter_out_expected[ 532] <= 18'h00000;
	 filter_out_expected[ 533] <= 18'h00000;
	 filter_out_expected[ 534] <= 18'h00000;
	 filter_out_expected[ 535] <= 18'h00000;
	 filter_out_expected[ 536] <= 18'h00000;
	 filter_out_expected[ 537] <= 18'h00000;
	 filter_out_expected[ 538] <= 18'h00000;
	 filter_out_expected[ 539] <= 18'h00000;
	 filter_out_expected[ 540] <= 18'h00000;
	 filter_out_expected[ 541] <= 18'h00000;
	 filter_out_expected[ 542] <= 18'h00000;
	 filter_out_expected[ 543] <= 18'h00000;
	 filter_out_expected[ 544] <= 18'h00000;
	 filter_out_expected[ 545] <= 18'h00000;
	 filter_out_expected[ 546] <= 18'h00000;
	 filter_out_expected[ 547] <= 18'h00000;
	 filter_out_expected[ 548] <= 18'h00000;
	 filter_out_expected[ 549] <= 18'h00000;
	 filter_out_expected[ 550] <= 18'h00000;
	 filter_out_expected[ 551] <= 18'h00000;
	 filter_out_expected[ 552] <= 18'h00000;
	 filter_out_expected[ 553] <= 18'h00000;
	 filter_out_expected[ 554] <= 18'h00000;
	 filter_out_expected[ 555] <= 18'h00000;
	 filter_out_expected[ 556] <= 18'h00000;
	 filter_out_expected[ 557] <= 18'h00000;
	 filter_out_expected[ 558] <= 18'h00000;
	 filter_out_expected[ 559] <= 18'h00000;
	 filter_out_expected[ 560] <= 18'h00000;
	 filter_out_expected[ 561] <= 18'h00000;
	 filter_out_expected[ 562] <= 18'h00000;
	 filter_out_expected[ 563] <= 18'h00000;
	 filter_out_expected[ 564] <= 18'h00000;
	 filter_out_expected[ 565] <= 18'h00000;
	 filter_out_expected[ 566] <= 18'h00000;
	 filter_out_expected[ 567] <= 18'h00000;
	 filter_out_expected[ 568] <= 18'h00000;
	 filter_out_expected[ 569] <= 18'h00000;
	 filter_out_expected[ 570] <= 18'h00000;
	 filter_out_expected[ 571] <= 18'h00000;
	 filter_out_expected[ 572] <= 18'h00000;
	 filter_out_expected[ 573] <= 18'h00000;
	 filter_out_expected[ 574] <= 18'h00000;
	 filter_out_expected[ 575] <= 18'h00000;
	 filter_out_expected[ 576] <= 18'h00000;
	 filter_out_expected[ 577] <= 18'h00000;
	 filter_out_expected[ 578] <= 18'h00000;
	 filter_out_expected[ 579] <= 18'h00000;
	 filter_out_expected[ 580] <= 18'h00000;
	 filter_out_expected[ 581] <= 18'h00000;
	 filter_out_expected[ 582] <= 18'h00000;
	 filter_out_expected[ 583] <= 18'h00000;
	 filter_out_expected[ 584] <= 18'h00000;
	 filter_out_expected[ 585] <= 18'h00000;
	 filter_out_expected[ 586] <= 18'h00000;
	 filter_out_expected[ 587] <= 18'h00000;
	 filter_out_expected[ 588] <= 18'h00000;
	 filter_out_expected[ 589] <= 18'h00000;
	 filter_out_expected[ 590] <= 18'h00000;
	 filter_out_expected[ 591] <= 18'h00000;
	 filter_out_expected[ 592] <= 18'h00000;
	 filter_out_expected[ 593] <= 18'h00000;
	 filter_out_expected[ 594] <= 18'h00000;
	 filter_out_expected[ 595] <= 18'h00000;
	 filter_out_expected[ 596] <= 18'h00000;
	 filter_out_expected[ 597] <= 18'h00000;
	 filter_out_expected[ 598] <= 18'h00000;
	 filter_out_expected[ 599] <= 18'h00000;
	 filter_out_expected[ 600] <= 18'h00000;
	 filter_out_expected[ 601] <= 18'h00000;
	 filter_out_expected[ 602] <= 18'h00000;
	 filter_out_expected[ 603] <= 18'h00000;
	 filter_out_expected[ 604] <= 18'h00000;
	 filter_out_expected[ 605] <= 18'h00000;
	 filter_out_expected[ 606] <= 18'h00000;
	 filter_out_expected[ 607] <= 18'h00000;
	 filter_out_expected[ 608] <= 18'h00000;
	 filter_out_expected[ 609] <= 18'h00000;
	 filter_out_expected[ 610] <= 18'h00000;
	 filter_out_expected[ 611] <= 18'h00000;
	 filter_out_expected[ 612] <= 18'h00000;
	 filter_out_expected[ 613] <= 18'h00000;
	 filter_out_expected[ 614] <= 18'h00000;
	 filter_out_expected[ 615] <= 18'h00000;
	 filter_out_expected[ 616] <= 18'h00000;
	 filter_out_expected[ 617] <= 18'h00000;
	 filter_out_expected[ 618] <= 18'h00000;
	 filter_out_expected[ 619] <= 18'h00000;
	 filter_out_expected[ 620] <= 18'h00000;
	 filter_out_expected[ 621] <= 18'h00000;
	 filter_out_expected[ 622] <= 18'h00000;
	 filter_out_expected[ 623] <= 18'h00000;
	 filter_out_expected[ 624] <= 18'h00000;
	 filter_out_expected[ 625] <= 18'h00000;
	 filter_out_expected[ 626] <= 18'h00000;
	 filter_out_expected[ 627] <= 18'h00000;
	 filter_out_expected[ 628] <= 18'h00000;
	 filter_out_expected[ 629] <= 18'h00000;
	 filter_out_expected[ 630] <= 18'h00000;
	 filter_out_expected[ 631] <= 18'h00000;
	 filter_out_expected[ 632] <= 18'h00000;
	 filter_out_expected[ 633] <= 18'h00000;
	 filter_out_expected[ 634] <= 18'h00000;
	 filter_out_expected[ 635] <= 18'h00000;
	 filter_out_expected[ 636] <= 18'h00000;
	 filter_out_expected[ 637] <= 18'h00000;
	 filter_out_expected[ 638] <= 18'h00000;
	 filter_out_expected[ 639] <= 18'h00000;
	 filter_out_expected[ 640] <= 18'h00000;
	 filter_out_expected[ 641] <= 18'h00000;
	 filter_out_expected[ 642] <= 18'h00000;
	 filter_out_expected[ 643] <= 18'h00000;
	 filter_out_expected[ 644] <= 18'h00000;
	 filter_out_expected[ 645] <= 18'h00000;
	 filter_out_expected[ 646] <= 18'h00000;
	 filter_out_expected[ 647] <= 18'h00000;
	 filter_out_expected[ 648] <= 18'h00000;
	 filter_out_expected[ 649] <= 18'h00000;
	 filter_out_expected[ 650] <= 18'h00000;
	 filter_out_expected[ 651] <= 18'h00000;
	 filter_out_expected[ 652] <= 18'h00000;
	 filter_out_expected[ 653] <= 18'h00000;
	 filter_out_expected[ 654] <= 18'h00000;
	 filter_out_expected[ 655] <= 18'h00000;
	 filter_out_expected[ 656] <= 18'h00000;
	 filter_out_expected[ 657] <= 18'h00000;
	 filter_out_expected[ 658] <= 18'h00000;
	 filter_out_expected[ 659] <= 18'h00000;
	 filter_out_expected[ 660] <= 18'h00000;
	 filter_out_expected[ 661] <= 18'h00000;
	 filter_out_expected[ 662] <= 18'h00000;
	 filter_out_expected[ 663] <= 18'h00000;
	 filter_out_expected[ 664] <= 18'h00000;
	 filter_out_expected[ 665] <= 18'h00000;
	 filter_out_expected[ 666] <= 18'h00000;
	 filter_out_expected[ 667] <= 18'h00000;
	 filter_out_expected[ 668] <= 18'h00000;
	 filter_out_expected[ 669] <= 18'h00000;
	 filter_out_expected[ 670] <= 18'h00000;
	 filter_out_expected[ 671] <= 18'h00000;
	 filter_out_expected[ 672] <= 18'h00000;
	 filter_out_expected[ 673] <= 18'h00000;
	 filter_out_expected[ 674] <= 18'h00000;
	 filter_out_expected[ 675] <= 18'h00000;
	 filter_out_expected[ 676] <= 18'h00000;
	 filter_out_expected[ 677] <= 18'h00000;
	 filter_out_expected[ 678] <= 18'h00000;
	 filter_out_expected[ 679] <= 18'h00000;
	 filter_out_expected[ 680] <= 18'h00000;
	 filter_out_expected[ 681] <= 18'h00000;
	 filter_out_expected[ 682] <= 18'h00000;
	 filter_out_expected[ 683] <= 18'h00000;
	 filter_out_expected[ 684] <= 18'h00000;
	 filter_out_expected[ 685] <= 18'h00000;
	 filter_out_expected[ 686] <= 18'h00000;
	 filter_out_expected[ 687] <= 18'h00000;
	 filter_out_expected[ 688] <= 18'h00000;
	 filter_out_expected[ 689] <= 18'h00000;
	 filter_out_expected[ 690] <= 18'h00000;
	 filter_out_expected[ 691] <= 18'h00000;
	 filter_out_expected[ 692] <= 18'h00000;
	 filter_out_expected[ 693] <= 18'h00000;
	 filter_out_expected[ 694] <= 18'h00000;
	 filter_out_expected[ 695] <= 18'h00000;
	 filter_out_expected[ 696] <= 18'h00000;
	 filter_out_expected[ 697] <= 18'h00000;
	 filter_out_expected[ 698] <= 18'h00000;
	 filter_out_expected[ 699] <= 18'h00000;
	 filter_out_expected[ 700] <= 18'h00000;
	 filter_out_expected[ 701] <= 18'h00000;
	 filter_out_expected[ 702] <= 18'h00000;
	 filter_out_expected[ 703] <= 18'h00000;
	 filter_out_expected[ 704] <= 18'h00000;
	 filter_out_expected[ 705] <= 18'h00000;
	 filter_out_expected[ 706] <= 18'h00000;
	 filter_out_expected[ 707] <= 18'h00000;
	 filter_out_expected[ 708] <= 18'h00000;
	 filter_out_expected[ 709] <= 18'h00000;
	 filter_out_expected[ 710] <= 18'h00000;
	 filter_out_expected[ 711] <= 18'h00000;
	 filter_out_expected[ 712] <= 18'h00000;
	 filter_out_expected[ 713] <= 18'h00000;
	 filter_out_expected[ 714] <= 18'h00000;
	 filter_out_expected[ 715] <= 18'h00000;
	 filter_out_expected[ 716] <= 18'h00000;
	 filter_out_expected[ 717] <= 18'h00000;
	 filter_out_expected[ 718] <= 18'h00000;
	 filter_out_expected[ 719] <= 18'h00000;
	 filter_out_expected[ 720] <= 18'h00000;
	 filter_out_expected[ 721] <= 18'h00000;
	 filter_out_expected[ 722] <= 18'h00000;
	 filter_out_expected[ 723] <= 18'h00000;
	 filter_out_expected[ 724] <= 18'h00000;
	 filter_out_expected[ 725] <= 18'h00000;
	 filter_out_expected[ 726] <= 18'h00000;
	 filter_out_expected[ 727] <= 18'h00000;
	 filter_out_expected[ 728] <= 18'h00000;
	 filter_out_expected[ 729] <= 18'h00000;
	 filter_out_expected[ 730] <= 18'h00000;
	 filter_out_expected[ 731] <= 18'h00000;
	 filter_out_expected[ 732] <= 18'h00000;
	 filter_out_expected[ 733] <= 18'h00000;
	 filter_out_expected[ 734] <= 18'h00000;
	 filter_out_expected[ 735] <= 18'h00000;
	 filter_out_expected[ 736] <= 18'h00000;
	 filter_out_expected[ 737] <= 18'h00000;
	 filter_out_expected[ 738] <= 18'h00000;
	 filter_out_expected[ 739] <= 18'h00000;
	 filter_out_expected[ 740] <= 18'h00000;
	 filter_out_expected[ 741] <= 18'h00000;
	 filter_out_expected[ 742] <= 18'h00000;
	 filter_out_expected[ 743] <= 18'h00000;
	 filter_out_expected[ 744] <= 18'h00000;
	 filter_out_expected[ 745] <= 18'h00000;
	 filter_out_expected[ 746] <= 18'h00000;
	 filter_out_expected[ 747] <= 18'h00000;
	 filter_out_expected[ 748] <= 18'h00000;
	 filter_out_expected[ 749] <= 18'h00000;
	 filter_out_expected[ 750] <= 18'h00000;
	 filter_out_expected[ 751] <= 18'h00000;
	 filter_out_expected[ 752] <= 18'h00000;
	 filter_out_expected[ 753] <= 18'h00000;
	 filter_out_expected[ 754] <= 18'h00000;
	 filter_out_expected[ 755] <= 18'h00000;
	 filter_out_expected[ 756] <= 18'h00000;
	 filter_out_expected[ 757] <= 18'h00000;
	 filter_out_expected[ 758] <= 18'h00000;
	 filter_out_expected[ 759] <= 18'h00000;
	 filter_out_expected[ 760] <= 18'h00000;
	 filter_out_expected[ 761] <= 18'h00000;
	 filter_out_expected[ 762] <= 18'h00000;
	 filter_out_expected[ 763] <= 18'h00000;
	 filter_out_expected[ 764] <= 18'h00000;
	 filter_out_expected[ 765] <= 18'h00000;
	 filter_out_expected[ 766] <= 18'h00000;
	 filter_out_expected[ 767] <= 18'h00000;
	 filter_out_expected[ 768] <= 18'h00000;
	 filter_out_expected[ 769] <= 18'h00000;
	 filter_out_expected[ 770] <= 18'h00000;
	 filter_out_expected[ 771] <= 18'h00000;
	 filter_out_expected[ 772] <= 18'h00000;
	 filter_out_expected[ 773] <= 18'h00000;
	 filter_out_expected[ 774] <= 18'h00000;
	 filter_out_expected[ 775] <= 18'h00000;
	 filter_out_expected[ 776] <= 18'h00000;
	 filter_out_expected[ 777] <= 18'h00000;
	 filter_out_expected[ 778] <= 18'h00000;
	 filter_out_expected[ 779] <= 18'h00000;
	 filter_out_expected[ 780] <= 18'h00000;
	 filter_out_expected[ 781] <= 18'h00000;
	 filter_out_expected[ 782] <= 18'h00000;
	 filter_out_expected[ 783] <= 18'h00000;
	 filter_out_expected[ 784] <= 18'h00000;
	 filter_out_expected[ 785] <= 18'h00000;
	 filter_out_expected[ 786] <= 18'h00000;
	 filter_out_expected[ 787] <= 18'h00000;
	 filter_out_expected[ 788] <= 18'h00000;
	 filter_out_expected[ 789] <= 18'h00000;
	 filter_out_expected[ 790] <= 18'h00000;
	 filter_out_expected[ 791] <= 18'h00000;
	 filter_out_expected[ 792] <= 18'h00000;
	 filter_out_expected[ 793] <= 18'h00000;
	 filter_out_expected[ 794] <= 18'h00000;
	 filter_out_expected[ 795] <= 18'h00000;
	 filter_out_expected[ 796] <= 18'h00000;
	 filter_out_expected[ 797] <= 18'h00000;
	 filter_out_expected[ 798] <= 18'h00000;
	 filter_out_expected[ 799] <= 18'h00000;
	 filter_out_expected[ 800] <= 18'h00000;
	 filter_out_expected[ 801] <= 18'h00000;
	 filter_out_expected[ 802] <= 18'h00000;
	 filter_out_expected[ 803] <= 18'h00000;
	 filter_out_expected[ 804] <= 18'h00000;
	 filter_out_expected[ 805] <= 18'h00000;
	 filter_out_expected[ 806] <= 18'h00000;
	 filter_out_expected[ 807] <= 18'h00000;
	 filter_out_expected[ 808] <= 18'h00000;
	 filter_out_expected[ 809] <= 18'h00000;
	 filter_out_expected[ 810] <= 18'h00000;
	 filter_out_expected[ 811] <= 18'h00000;
	 filter_out_expected[ 812] <= 18'h00000;
	 filter_out_expected[ 813] <= 18'h00000;
	 filter_out_expected[ 814] <= 18'h00000;
	 filter_out_expected[ 815] <= 18'h00000;
	 filter_out_expected[ 816] <= 18'h00000;
	 filter_out_expected[ 817] <= 18'h00000;
	 filter_out_expected[ 818] <= 18'h00000;
	 filter_out_expected[ 819] <= 18'h00000;
	 filter_out_expected[ 820] <= 18'h00000;
	 filter_out_expected[ 821] <= 18'h00000;
	 filter_out_expected[ 822] <= 18'h00000;
	 filter_out_expected[ 823] <= 18'h00000;
	 filter_out_expected[ 824] <= 18'h00000;
	 filter_out_expected[ 825] <= 18'h00000;
	 filter_out_expected[ 826] <= 18'h00000;
	 filter_out_expected[ 827] <= 18'h00000;
	 filter_out_expected[ 828] <= 18'h00000;
	 filter_out_expected[ 829] <= 18'h00000;
	 filter_out_expected[ 830] <= 18'h00000;
	 filter_out_expected[ 831] <= 18'h00000;
	 filter_out_expected[ 832] <= 18'h00000;
	 filter_out_expected[ 833] <= 18'h00000;
	 filter_out_expected[ 834] <= 18'h00000;
	 filter_out_expected[ 835] <= 18'h00000;
	 filter_out_expected[ 836] <= 18'h00000;
	 filter_out_expected[ 837] <= 18'h00000;
	 filter_out_expected[ 838] <= 18'h00000;
	 filter_out_expected[ 839] <= 18'h00000;
	 filter_out_expected[ 840] <= 18'h00000;
	 filter_out_expected[ 841] <= 18'h00000;
	 filter_out_expected[ 842] <= 18'h00000;
	 filter_out_expected[ 843] <= 18'h00000;
	 filter_out_expected[ 844] <= 18'h00000;
	 filter_out_expected[ 845] <= 18'h00000;
	 filter_out_expected[ 846] <= 18'h00000;
	 filter_out_expected[ 847] <= 18'h00000;
	 filter_out_expected[ 848] <= 18'h00000;
	 filter_out_expected[ 849] <= 18'h00000;
	 filter_out_expected[ 850] <= 18'h00000;
	 filter_out_expected[ 851] <= 18'h00000;
	 filter_out_expected[ 852] <= 18'h00000;
	 filter_out_expected[ 853] <= 18'h00000;
	 filter_out_expected[ 854] <= 18'h00000;
	 filter_out_expected[ 855] <= 18'h00000;
	 filter_out_expected[ 856] <= 18'h00000;
	 filter_out_expected[ 857] <= 18'h00000;
	 filter_out_expected[ 858] <= 18'h00000;
	 filter_out_expected[ 859] <= 18'h00000;
	 filter_out_expected[ 860] <= 18'h00000;
	 filter_out_expected[ 861] <= 18'h00000;
	 filter_out_expected[ 862] <= 18'h00000;
	 filter_out_expected[ 863] <= 18'h00000;
	 filter_out_expected[ 864] <= 18'h00000;
	 filter_out_expected[ 865] <= 18'h00000;
	 filter_out_expected[ 866] <= 18'h00000;
	 filter_out_expected[ 867] <= 18'h00000;
	 filter_out_expected[ 868] <= 18'h00000;
	 filter_out_expected[ 869] <= 18'h00000;
	 filter_out_expected[ 870] <= 18'h00000;
	 filter_out_expected[ 871] <= 18'h00000;
	 filter_out_expected[ 872] <= 18'h00000;
	 filter_out_expected[ 873] <= 18'h00000;
	 filter_out_expected[ 874] <= 18'h00000;
	 filter_out_expected[ 875] <= 18'h00000;
	 filter_out_expected[ 876] <= 18'h00000;
	 filter_out_expected[ 877] <= 18'h00000;
	 filter_out_expected[ 878] <= 18'h00000;
	 filter_out_expected[ 879] <= 18'h00000;
	 filter_out_expected[ 880] <= 18'h00000;
	 filter_out_expected[ 881] <= 18'h00000;
	 filter_out_expected[ 882] <= 18'h00000;
	 filter_out_expected[ 883] <= 18'h00000;
	 filter_out_expected[ 884] <= 18'h00000;
	 filter_out_expected[ 885] <= 18'h00000;
	 filter_out_expected[ 886] <= 18'h00000;
	 filter_out_expected[ 887] <= 18'h00000;
	 filter_out_expected[ 888] <= 18'h00000;
	 filter_out_expected[ 889] <= 18'h00000;
	 filter_out_expected[ 890] <= 18'h00000;
	 filter_out_expected[ 891] <= 18'h00000;
	 filter_out_expected[ 892] <= 18'h00000;
	 filter_out_expected[ 893] <= 18'h00000;
	 filter_out_expected[ 894] <= 18'h00000;
	 filter_out_expected[ 895] <= 18'h00000;
	 filter_out_expected[ 896] <= 18'h00000;
	 filter_out_expected[ 897] <= 18'h00000;
	 filter_out_expected[ 898] <= 18'h00000;
	 filter_out_expected[ 899] <= 18'h00000;
	 filter_out_expected[ 900] <= 18'h00000;
	 filter_out_expected[ 901] <= 18'h00000;
	 filter_out_expected[ 902] <= 18'h00000;
	 filter_out_expected[ 903] <= 18'h00000;
	 filter_out_expected[ 904] <= 18'h00000;
	 filter_out_expected[ 905] <= 18'h00000;
	 filter_out_expected[ 906] <= 18'h00000;
	 filter_out_expected[ 907] <= 18'h00000;
	 filter_out_expected[ 908] <= 18'h00000;
	 filter_out_expected[ 909] <= 18'h00000;
	 filter_out_expected[ 910] <= 18'h00000;
	 filter_out_expected[ 911] <= 18'h00000;
	 filter_out_expected[ 912] <= 18'h00000;
	 filter_out_expected[ 913] <= 18'h00000;
	 filter_out_expected[ 914] <= 18'h00000;
	 filter_out_expected[ 915] <= 18'h00000;
	 filter_out_expected[ 916] <= 18'h00000;
	 filter_out_expected[ 917] <= 18'h00000;
	 filter_out_expected[ 918] <= 18'h00000;
	 filter_out_expected[ 919] <= 18'h00000;
	 filter_out_expected[ 920] <= 18'h00000;
	 filter_out_expected[ 921] <= 18'h00000;
	 filter_out_expected[ 922] <= 18'h00000;
	 filter_out_expected[ 923] <= 18'h00000;
	 filter_out_expected[ 924] <= 18'h00000;
	 filter_out_expected[ 925] <= 18'h00000;
	 filter_out_expected[ 926] <= 18'h00000;
	 filter_out_expected[ 927] <= 18'h00000;
	 filter_out_expected[ 928] <= 18'h00000;
	 filter_out_expected[ 929] <= 18'h00000;
	 filter_out_expected[ 930] <= 18'h00000;
	 filter_out_expected[ 931] <= 18'h00000;
	 filter_out_expected[ 932] <= 18'h00000;
	 filter_out_expected[ 933] <= 18'h00000;
	 filter_out_expected[ 934] <= 18'h00000;
	 filter_out_expected[ 935] <= 18'h00000;
	 filter_out_expected[ 936] <= 18'h00000;
	 filter_out_expected[ 937] <= 18'h00000;
	 filter_out_expected[ 938] <= 18'h00000;
	 filter_out_expected[ 939] <= 18'h00000;
	 filter_out_expected[ 940] <= 18'h00000;
	 filter_out_expected[ 941] <= 18'h00000;
	 filter_out_expected[ 942] <= 18'h00000;
	 filter_out_expected[ 943] <= 18'h00000;
	 filter_out_expected[ 944] <= 18'h00000;
	 filter_out_expected[ 945] <= 18'h00000;
	 filter_out_expected[ 946] <= 18'h00000;
	 filter_out_expected[ 947] <= 18'h00000;
	 filter_out_expected[ 948] <= 18'h00000;
	 filter_out_expected[ 949] <= 18'h00000;
	 filter_out_expected[ 950] <= 18'h00000;
	 filter_out_expected[ 951] <= 18'h00000;
	 filter_out_expected[ 952] <= 18'h00000;
	 filter_out_expected[ 953] <= 18'h00000;
	 filter_out_expected[ 954] <= 18'h00000;
	 filter_out_expected[ 955] <= 18'h00000;
	 filter_out_expected[ 956] <= 18'h00000;
	 filter_out_expected[ 957] <= 18'h00000;
	 filter_out_expected[ 958] <= 18'h00000;
	 filter_out_expected[ 959] <= 18'h00000;
	 filter_out_expected[ 960] <= 18'h00000;
	 filter_out_expected[ 961] <= 18'h00000;
	 filter_out_expected[ 962] <= 18'h00000;
	 filter_out_expected[ 963] <= 18'h00000;
	 filter_out_expected[ 964] <= 18'h00000;
	 filter_out_expected[ 965] <= 18'h00000;
	 filter_out_expected[ 966] <= 18'h00000;
	 filter_out_expected[ 967] <= 18'h00000;
	 filter_out_expected[ 968] <= 18'h00000;
	 filter_out_expected[ 969] <= 18'h00000;
	 filter_out_expected[ 970] <= 18'h00000;
	 filter_out_expected[ 971] <= 18'h00000;
	 filter_out_expected[ 972] <= 18'h00000;
	 filter_out_expected[ 973] <= 18'h00000;
	 filter_out_expected[ 974] <= 18'h00000;
	 filter_out_expected[ 975] <= 18'h00000;
	 filter_out_expected[ 976] <= 18'h00000;
	 filter_out_expected[ 977] <= 18'h00000;
	 filter_out_expected[ 978] <= 18'h00000;
	 filter_out_expected[ 979] <= 18'h00000;
	 filter_out_expected[ 980] <= 18'h00000;
	 filter_out_expected[ 981] <= 18'h00000;
	 filter_out_expected[ 982] <= 18'h00000;
	 filter_out_expected[ 983] <= 18'h00000;
	 filter_out_expected[ 984] <= 18'h00000;
	 filter_out_expected[ 985] <= 18'h00000;
	 filter_out_expected[ 986] <= 18'h00000;
	 filter_out_expected[ 987] <= 18'h00000;
	 filter_out_expected[ 988] <= 18'h00000;
	 filter_out_expected[ 989] <= 18'h00000;
	 filter_out_expected[ 990] <= 18'h00000;
	 filter_out_expected[ 991] <= 18'h00000;
	 filter_out_expected[ 992] <= 18'h00000;
	 filter_out_expected[ 993] <= 18'h00000;
	 filter_out_expected[ 994] <= 18'h00000;
	 filter_out_expected[ 995] <= 18'h00000;
	 filter_out_expected[ 996] <= 18'h00000;
	 filter_out_expected[ 997] <= 18'h00000;
	 filter_out_expected[ 998] <= 18'h00000;
	 filter_out_expected[ 999] <= 18'h00000;
	 filter_out_expected[1000] <= 18'h00000;
	 filter_out_expected[1001] <= 18'h00000;
	 filter_out_expected[1002] <= 18'h00000;
	 filter_out_expected[1003] <= 18'h00000;
	 filter_out_expected[1004] <= 18'h00000;
	 filter_out_expected[1005] <= 18'h00000;
	 filter_out_expected[1006] <= 18'h00000;
	 filter_out_expected[1007] <= 18'h00000;
	 filter_out_expected[1008] <= 18'h00000;
	 filter_out_expected[1009] <= 18'h00000;
	 filter_out_expected[1010] <= 18'h00000;
	 filter_out_expected[1011] <= 18'h00000;
	 filter_out_expected[1012] <= 18'h00000;
	 filter_out_expected[1013] <= 18'h00000;
	 filter_out_expected[1014] <= 18'h00000;
	 filter_out_expected[1015] <= 18'h00000;
	 filter_out_expected[1016] <= 18'h00000;
	 filter_out_expected[1017] <= 18'h00000;
	 filter_out_expected[1018] <= 18'h00000;
	 filter_out_expected[1019] <= 18'h00000;
	 filter_out_expected[1020] <= 18'h00000;
	 filter_out_expected[1021] <= 18'h00000;
	 filter_out_expected[1022] <= 18'h00000;
	 filter_out_expected[1023] <= 18'h00000;
	 filter_out_expected[1024] <= 18'h00000;
	 filter_out_expected[1025] <= 18'h00000;
	 filter_out_expected[1026] <= 18'h00000;
	 filter_out_expected[1027] <= 18'h00000;
	 filter_out_expected[1028] <= 18'h00000;
	 filter_out_expected[1029] <= 18'h00000;
	 filter_out_expected[1030] <= 18'h00000;
	 filter_out_expected[1031] <= 18'h00000;
	 filter_out_expected[1032] <= 18'h00000;
	 filter_out_expected[1033] <= 18'h00000;
	 filter_out_expected[1034] <= 18'h00000;
	 filter_out_expected[1035] <= 18'h00000;
	 filter_out_expected[1036] <= 18'h00000;
	 filter_out_expected[1037] <= 18'h00000;
	 filter_out_expected[1038] <= 18'h00000;
	 filter_out_expected[1039] <= 18'h00000;
	 filter_out_expected[1040] <= 18'h00000;
	 filter_out_expected[1041] <= 18'h00000;
	 filter_out_expected[1042] <= 18'h00000;
	 filter_out_expected[1043] <= 18'h00000;
	 filter_out_expected[1044] <= 18'h00000;
	 filter_out_expected[1045] <= 18'h00000;
	 filter_out_expected[1046] <= 18'h00000;
	 filter_out_expected[1047] <= 18'h00000;
	 filter_out_expected[1048] <= 18'h00000;
	 filter_out_expected[1049] <= 18'h00000;
	 filter_out_expected[1050] <= 18'h00000;
	 filter_out_expected[1051] <= 18'h00000;
	 filter_out_expected[1052] <= 18'h00000;
	 filter_out_expected[1053] <= 18'h00000;
	 filter_out_expected[1054] <= 18'h00000;
	 filter_out_expected[1055] <= 18'h00000;
	 filter_out_expected[1056] <= 18'h00000;
	 filter_out_expected[1057] <= 18'h00000;
	 filter_out_expected[1058] <= 18'h00000;
	 filter_out_expected[1059] <= 18'h00000;
	 filter_out_expected[1060] <= 18'h00000;
	 filter_out_expected[1061] <= 18'h00000;
	 filter_out_expected[1062] <= 18'h00000;
	 filter_out_expected[1063] <= 18'h00000;
	 filter_out_expected[1064] <= 18'h00000;
	 filter_out_expected[1065] <= 18'h00000;
	 filter_out_expected[1066] <= 18'h00000;
	 filter_out_expected[1067] <= 18'h00000;
	 filter_out_expected[1068] <= 18'h03018;
	 filter_out_expected[1069] <= 18'h0b070;
	 filter_out_expected[1070] <= 18'h13108;
	 filter_out_expected[1071] <= 18'h131a0;
	 filter_out_expected[1072] <= 18'h081e0;
	 filter_out_expected[1073] <= 18'h381a0;
	 filter_out_expected[1074] <= 18'h2d108;
	 filter_out_expected[1075] <= 18'h2d070;
	 filter_out_expected[1076] <= 18'h35018;
	 filter_out_expected[1077] <= 18'h3d000;
	 filter_out_expected[1078] <= 18'h00000;
	 filter_out_expected[1079] <= 18'h3d000;
	 filter_out_expected[1080] <= 18'h35000;
	 filter_out_expected[1081] <= 18'h2d001;
	 filter_out_expected[1082] <= 18'h2d002;
	 filter_out_expected[1083] <= 18'h38007;
	 filter_out_expected[1084] <= 18'h08014;
	 filter_out_expected[1085] <= 18'h13031;
	 filter_out_expected[1086] <= 18'h13063;
	 filter_out_expected[1087] <= 18'h0b0ae;
	 filter_out_expected[1088] <= 18'h03115;
	 filter_out_expected[1089] <= 18'h00199;
	 filter_out_expected[1090] <= 18'h0023a;
	 filter_out_expected[1091] <= 18'h002f7;
	 filter_out_expected[1092] <= 18'h003d1;
	 filter_out_expected[1093] <= 18'h004c6;
	 filter_out_expected[1094] <= 18'h005d5;
	 filter_out_expected[1095] <= 18'h006fc;
	 filter_out_expected[1096] <= 18'h0083b;
	 filter_out_expected[1097] <= 18'h0098e;
	 filter_out_expected[1098] <= 18'h00af3;
	 filter_out_expected[1099] <= 18'h00c65;
	 filter_out_expected[1100] <= 18'h00de0;
	 filter_out_expected[1101] <= 18'h00f5f;
	 filter_out_expected[1102] <= 18'h010da;
	 filter_out_expected[1103] <= 18'h0124a;
	 filter_out_expected[1104] <= 18'h013a7;
	 filter_out_expected[1105] <= 18'h014e7;
	 filter_out_expected[1106] <= 18'h015fe;
	 filter_out_expected[1107] <= 18'h016e1;
	 filter_out_expected[1108] <= 18'h01784;
	 filter_out_expected[1109] <= 18'h017d7;
	 filter_out_expected[1110] <= 18'h017ce;
	 filter_out_expected[1111] <= 18'h01759;
	 filter_out_expected[1112] <= 18'h0166a;
	 filter_out_expected[1113] <= 18'h014f2;
	 filter_out_expected[1114] <= 18'h012e5;
	 filter_out_expected[1115] <= 18'h01036;
	 filter_out_expected[1116] <= 18'h00cdd;
	 filter_out_expected[1117] <= 18'h008d2;
	 filter_out_expected[1118] <= 18'h00413;
	 filter_out_expected[1119] <= 18'h3fea2;
	 filter_out_expected[1120] <= 18'h3f886;
	 filter_out_expected[1121] <= 18'h3f1cc;
	 filter_out_expected[1122] <= 18'h3ea88;
	 filter_out_expected[1123] <= 18'h3e2d6;
	 filter_out_expected[1124] <= 18'h3dada;
	 filter_out_expected[1125] <= 18'h3d2c1;
	 filter_out_expected[1126] <= 18'h3cabf;
	 filter_out_expected[1127] <= 18'h3c311;
	 filter_out_expected[1128] <= 18'h3bbfa;
	 filter_out_expected[1129] <= 18'h3b5c3;
	 filter_out_expected[1130] <= 18'h3b0bb;
	 filter_out_expected[1131] <= 18'h3ad33;
	 filter_out_expected[1132] <= 18'h3ab79;
	 filter_out_expected[1133] <= 18'h3abd8;
	 filter_out_expected[1134] <= 18'h3ae93;
	 filter_out_expected[1135] <= 18'h3b3e2;
	 filter_out_expected[1136] <= 18'h3bbe9;
	 filter_out_expected[1137] <= 18'h3c6bb;
	 filter_out_expected[1138] <= 18'h3d450;
	 filter_out_expected[1139] <= 18'h3e481;
	 filter_out_expected[1140] <= 18'h3f707;
	 filter_out_expected[1141] <= 18'h00b7a;
	 filter_out_expected[1142] <= 18'h0214a;
	 filter_out_expected[1143] <= 18'h037c6;
	 filter_out_expected[1144] <= 18'h04e1d;
	 filter_out_expected[1145] <= 18'h06360;
	 filter_out_expected[1146] <= 18'h07690;
	 filter_out_expected[1147] <= 18'h0869f;
	 filter_out_expected[1148] <= 18'h09285;
	 filter_out_expected[1149] <= 18'h09949;
	 filter_out_expected[1150] <= 18'h09a12;
	 filter_out_expected[1151] <= 18'h09439;
	 filter_out_expected[1152] <= 18'h08759;
	 filter_out_expected[1153] <= 18'h0735e;
	 filter_out_expected[1154] <= 18'h05892;
	 filter_out_expected[1155] <= 18'h037ab;
	 filter_out_expected[1156] <= 18'h011c8;
	 filter_out_expected[1157] <= 18'h3e875;
	 filter_out_expected[1158] <= 18'h3bda2;
	 filter_out_expected[1159] <= 18'h3938d;
	 filter_out_expected[1160] <= 18'h36cac;
	 filter_out_expected[1161] <= 18'h34b8e;
	 filter_out_expected[1162] <= 18'h332ad;
	 filter_out_expected[1163] <= 18'h32443;
	 filter_out_expected[1164] <= 18'h3221c;
	 filter_out_expected[1165] <= 18'h32d67;
	 filter_out_expected[1166] <= 18'h34689;
	 filter_out_expected[1167] <= 18'h36cfd;
	 filter_out_expected[1168] <= 18'h39f41;
	 filter_out_expected[1169] <= 18'h3dad0;
	 filter_out_expected[1170] <= 18'h01c34;
	 filter_out_expected[1171] <= 18'h05f31;
	 filter_out_expected[1172] <= 18'h09efa;
	 filter_out_expected[1173] <= 18'h0d689;
	 filter_out_expected[1174] <= 18'h10101;
	 filter_out_expected[1175] <= 18'h11a17;
	 filter_out_expected[1176] <= 18'h11e85;
	 filter_out_expected[1177] <= 18'h10c6e;
	 filter_out_expected[1178] <= 18'h0e3b1;
	 filter_out_expected[1179] <= 18'h0a624;
	 filter_out_expected[1180] <= 18'h0579a;
	 filter_out_expected[1181] <= 18'h3fdc8;
	 filter_out_expected[1182] <= 18'h39fee;
	 filter_out_expected[1183] <= 18'h34651;
	 filter_out_expected[1184] <= 18'h2f989;
	 filter_out_expected[1185] <= 18'h2c1b0;
	 filter_out_expected[1186] <= 18'h2a583;
	 filter_out_expected[1187] <= 18'h2a98f;
	 filter_out_expected[1188] <= 18'h2cf7a;
	 filter_out_expected[1189] <= 18'h3158d;
	 filter_out_expected[1190] <= 18'h37689;
	 filter_out_expected[1191] <= 18'h3e9e3;
	 filter_out_expected[1192] <= 18'h0645c;
	 filter_out_expected[1193] <= 18'h0d909;
	 filter_out_expected[1194] <= 18'h13aa0;
	 filter_out_expected[1195] <= 18'h17cff;
	 filter_out_expected[1196] <= 18'h196b7;
	 filter_out_expected[1197] <= 18'h1826f;
	 filter_out_expected[1198] <= 18'h13ff2;
	 filter_out_expected[1199] <= 18'h0d4ac;
	 filter_out_expected[1200] <= 18'h04b80;
	 filter_out_expected[1201] <= 18'h3b3e6;
	 filter_out_expected[1202] <= 18'h3204a;
	 filter_out_expected[1203] <= 18'h2a3e9;
	 filter_out_expected[1204] <= 18'h25048;
	 filter_out_expected[1205] <= 18'h232ac;
	 filter_out_expected[1206] <= 18'h251e7;
	 filter_out_expected[1207] <= 18'h2acd4;
	 filter_out_expected[1208] <= 18'h339d2;
	 filter_out_expected[1209] <= 18'h3e773;
	 filter_out_expected[1210] <= 18'h09e64;
	 filter_out_expected[1211] <= 18'h14467;
	 filter_out_expected[1212] <= 18'h1c00f;
	 filter_out_expected[1213] <= 18'h1fcb5;
	 filter_out_expected[1214] <= 18'h1ee13;
	 filter_out_expected[1215] <= 18'h192da;
	 filter_out_expected[1216] <= 18'h0f5c9;
	 filter_out_expected[1217] <= 18'h02ce0;
	 filter_out_expected[1218] <= 18'h3569f;
	 filter_out_expected[1219] <= 18'h29596;
	 filter_out_expected[1220] <= 18'h20ae1;
	 filter_out_expected[1221] <= 18'h1d059;
	 filter_out_expected[1222] <= 18'h1f38e;
	 filter_out_expected[1223] <= 18'h2727b;
	 filter_out_expected[1224] <= 18'h33abc;
	 filter_out_expected[1225] <= 18'h02bb2;
	 filter_out_expected[1226] <= 18'h11b79;
	 filter_out_expected[1227] <= 18'h1de03;
	 filter_out_expected[1228] <= 18'h24d43;
	 filter_out_expected[1229] <= 18'h250d3;
	 filter_out_expected[1230] <= 18'h1e3a5;
	 filter_out_expected[1231] <= 18'h1164f;
	 filter_out_expected[1232] <= 18'h00d42;
	 filter_out_expected[1233] <= 18'h2facb;
	 filter_out_expected[1234] <= 18'h215ca;
	 filter_out_expected[1235] <= 18'h18eb1;
	 filter_out_expected[1236] <= 18'h184fd;
	 filter_out_expected[1237] <= 18'h1ff78;
	 filter_out_expected[1238] <= 18'h2e926;
	 filter_out_expected[1239] <= 18'h0140c;
	 filter_out_expected[1240] <= 18'h141a9;
	 filter_out_expected[1241] <= 18'h22fc7;
	 filter_out_expected[1242] <= 18'h2a71e;
	 filter_out_expected[1243] <= 18'h2888b;
	 filter_out_expected[1244] <= 18'h1d5bd;
	 filter_out_expected[1245] <= 18'h0b2c8;
	 filter_out_expected[1246] <= 18'h35fc2;
	 filter_out_expected[1247] <= 18'h22b2a;
	 filter_out_expected[1248] <= 18'h15fdb;
	 filter_out_expected[1249] <= 18'h13294;
	 filter_out_expected[1250] <= 18'h1b3b0;
	 filter_out_expected[1251] <= 18'h2c8ef;
	 filter_out_expected[1252] <= 18'h031ab;
	 filter_out_expected[1253] <= 18'h19520;
	 filter_out_expected[1254] <= 18'h297fc;
	 filter_out_expected[1255] <= 18'h2f40d;
	 filter_out_expected[1256] <= 18'h28bf1;
	 filter_out_expected[1257] <= 18'h17531;
	 filter_out_expected[1258] <= 18'h3f535;
	 filter_out_expected[1259] <= 18'h270ef;
	 filter_out_expected[1260] <= 18'h152b8;
	 filter_out_expected[1261] <= 18'h0ecf6;
	 filter_out_expected[1262] <= 18'h1619f;
	 filter_out_expected[1263] <= 18'h29605;
	 filter_out_expected[1264] <= 18'h03761;
	 filter_out_expected[1265] <= 18'h1cffe;
	 filter_out_expected[1266] <= 18'h2e810;
	 filter_out_expected[1267] <= 18'h3292b;
	 filter_out_expected[1268] <= 18'h279e4;
	 filter_out_expected[1269] <= 18'h1088e;
	 filter_out_expected[1270] <= 18'h34093;
	 filter_out_expected[1271] <= 18'h1ac34;
	 filter_out_expected[1272] <= 18'h0cac3;
	 filter_out_expected[1273] <= 18'h0e7ea;
	 filter_out_expected[1274] <= 18'h20108;
	 filter_out_expected[1275] <= 18'h3c257;
	 filter_out_expected[1276] <= 18'h19e62;
	 filter_out_expected[1277] <= 18'h2f9dd;
	 filter_out_expected[1278] <= 18'h35e93;
	 filter_out_expected[1279] <= 18'h2a4bf;
	 filter_out_expected[1280] <= 18'h10417;
	 filter_out_expected[1281] <= 18'h30506;
	 filter_out_expected[1282] <= 18'h15533;
	 filter_out_expected[1283] <= 18'h08c91;
	 filter_out_expected[1284] <= 18'h0f6f5;
	 filter_out_expected[1285] <= 18'h275ce;
	 filter_out_expected[1286] <= 18'h08682;
	 filter_out_expected[1287] <= 18'h26d79;
	 filter_out_expected[1288] <= 18'h3783f;
	 filter_out_expected[1289] <= 18'h33fc5;
	 filter_out_expected[1290] <= 18'h1d1ec;
	 filter_out_expected[1291] <= 18'h3b120;
	 filter_out_expected[1292] <= 18'h1a7ae;
	 filter_out_expected[1293] <= 18'h07d34;
	 filter_out_expected[1294] <= 18'h0a96b;
	 filter_out_expected[1295] <= 18'h2223e;
	 filter_out_expected[1296] <= 18'h05a9f;
	 filter_out_expected[1297] <= 18'h2755d;
	 filter_out_expected[1298] <= 18'h39a99;
	 filter_out_expected[1299] <= 18'h34f3c;
	 filter_out_expected[1300] <= 18'h1aab2;
	 filter_out_expected[1301] <= 18'h352df;
	 filter_out_expected[1302] <= 18'h13ca8;
	 filter_out_expected[1303] <= 18'h04866;
	 filter_out_expected[1304] <= 18'h0e26f;
	 filter_out_expected[1305] <= 18'h2d0a9;
	 filter_out_expected[1306] <= 18'h14573;
	 filter_out_expected[1307] <= 18'h3335e;
	 filter_out_expected[1308] <= 18'h3c0a3;
	 filter_out_expected[1309] <= 18'h2a8ed;
	 filter_out_expected[1310] <= 18'h060f7;
	 filter_out_expected[1311] <= 18'h1e8b9;
	 filter_out_expected[1312] <= 18'h05c8b;
	 filter_out_expected[1313] <= 18'h07490;
	 filter_out_expected[1314] <= 18'h22cb6;
	 filter_out_expected[1315] <= 18'h0c040;
	 filter_out_expected[1316] <= 18'h2ff36;
	 filter_out_expected[1317] <= 18'h3d9fc;
	 filter_out_expected[1318] <= 18'h2e34d;
	 filter_out_expected[1319] <= 18'h089d3;
	 filter_out_expected[1320] <= 18'h1e9d4;
	 filter_out_expected[1321] <= 18'h04887;
	 filter_out_expected[1322] <= 18'h075f2;
	 filter_out_expected[1323] <= 18'h26275;
	 filter_out_expected[1324] <= 18'h11f9a;
	 filter_out_expected[1325] <= 18'h350ef;
	 filter_out_expected[1326] <= 18'h3d8ee;
	 filter_out_expected[1327] <= 18'h26c75;
	 filter_out_expected[1328] <= 18'h3bfb6;
	 filter_out_expected[1329] <= 18'h13078;
	 filter_out_expected[1330] <= 18'h01492;
	 filter_out_expected[1331] <= 18'h105f1;
	 filter_out_expected[1332] <= 18'h38b9a;
	 filter_out_expected[1333] <= 18'h25267;
	 filter_out_expected[1334] <= 18'h3dd44;
	 filter_out_expected[1335] <= 18'h35294;
	 filter_out_expected[1336] <= 18'h0f78b;
	 filter_out_expected[1337] <= 18'h21206;
	 filter_out_expected[1338] <= 18'h03aea;
	 filter_out_expected[1339] <= 18'h07c12;
	 filter_out_expected[1340] <= 18'h2b6f0;
	 filter_out_expected[1341] <= 18'h1ae01;
	 filter_out_expected[1342] <= 18'h3b288;
	 filter_out_expected[1343] <= 18'h39943;
	 filter_out_expected[1344] <= 18'h16b1d;
	 filter_out_expected[1345] <= 18'h267d3;
	 filter_out_expected[1346] <= 18'h051ea;
	 filter_out_expected[1347] <= 18'h0675e;
	 filter_out_expected[1348] <= 18'h2a0d5;
	 filter_out_expected[1349] <= 18'h1ae18;
	 filter_out_expected[1350] <= 18'h3b95d;
	 filter_out_expected[1351] <= 18'h3820a;
	 filter_out_expected[1352] <= 18'h124cb;
	 filter_out_expected[1353] <= 18'h21206;
	 filter_out_expected[1354] <= 18'h030c3;
	 filter_out_expected[1355] <= 18'h0b08b;
	 filter_out_expected[1356] <= 18'h345f3;
	 filter_out_expected[1357] <= 18'h251f7;
	 filter_out_expected[1358] <= 18'h3e39b;
	 filter_out_expected[1359] <= 18'h2f5ce;
	 filter_out_expected[1360] <= 18'h01d9e;
	 filter_out_expected[1361] <= 18'h131d5;
	 filter_out_expected[1362] <= 18'h01cc3;
	 filter_out_expected[1363] <= 18'h198a6;
	 filter_out_expected[1364] <= 18'h0ad75;
	 filter_out_expected[1365] <= 18'h34e14;
	 filter_out_expected[1366] <= 18'h3b4b0;
	 filter_out_expected[1367] <= 18'h19824;
	 filter_out_expected[1368] <= 18'h26571;
	 filter_out_expected[1369] <= 18'h04d62;
	 filter_out_expected[1370] <= 18'h0c442;
	 filter_out_expected[1371] <= 18'h37af8;
	 filter_out_expected[1372] <= 18'h28dfb;
	 filter_out_expected[1373] <= 18'h3d2ea;
	 filter_out_expected[1374] <= 18'h260e6;
	 filter_out_expected[1375] <= 18'h33cca;
	 filter_out_expected[1376] <= 18'h0a670;
	 filter_out_expected[1377] <= 18'h07d80;
	 filter_out_expected[1378] <= 18'h2e272;
	 filter_out_expected[1379] <= 18'h21711;
	 filter_out_expected[1380] <= 18'h3bf67;
	 filter_out_expected[1381] <= 18'h29f45;
	 filter_out_expected[1382] <= 18'h38b1f;
	 filter_out_expected[1383] <= 18'h0d104;
	 filter_out_expected[1384] <= 18'h080a9;
	 filter_out_expected[1385] <= 18'h2d906;
	 filter_out_expected[1386] <= 18'h210eb;
	 filter_out_expected[1387] <= 18'h3aefc;
	 filter_out_expected[1388] <= 18'h271a1;
	 filter_out_expected[1389] <= 18'h34e4d;
	 filter_out_expected[1390] <= 18'h0b964;
	 filter_out_expected[1391] <= 18'h0bc29;
	 filter_out_expected[1392] <= 18'h355a1;
	 filter_out_expected[1393] <= 18'h27406;
	 filter_out_expected[1394] <= 18'h396db;
	 filter_out_expected[1395] <= 18'h1d2b1;
	 filter_out_expected[1396] <= 18'h295db;
	 filter_out_expected[1397] <= 18'h084f5;
	 filter_out_expected[1398] <= 18'h152bf;
	 filter_out_expected[1399] <= 18'h0559b;
	 filter_out_expected[1400] <= 18'h30d10;
	 filter_out_expected[1401] <= 18'h333bb;
	 filter_out_expected[1402] <= 18'h0a90d;
	 filter_out_expected[1403] <= 18'h19356;
	 filter_out_expected[1404] <= 18'h09240;
	 filter_out_expected[1405] <= 18'h2816e;
	 filter_out_expected[1406] <= 18'h1b673;
	 filter_out_expected[1407] <= 18'h36ad0;
	 filter_out_expected[1408] <= 18'h2234e;
	 filter_out_expected[1409] <= 18'h2ff56;
	 filter_out_expected[1410] <= 18'h0c2d2;
	 filter_out_expected[1411] <= 18'h167dd;
	 filter_out_expected[1412] <= 18'h05a62;
	 filter_out_expected[1413] <= 18'h2f65f;
	 filter_out_expected[1414] <= 18'h2e337;
	 filter_out_expected[1415] <= 18'h033cb;
	 filter_out_expected[1416] <= 18'h15acd;
	 filter_out_expected[1417] <= 18'h0f2d6;
	 filter_out_expected[1418] <= 18'h359b8;
	 filter_out_expected[1419] <= 18'h25507;
	 filter_out_expected[1420] <= 18'h31f09;
	 filter_out_expected[1421] <= 18'h0fce6;
	 filter_out_expected[1422] <= 18'h1f22e;
	 filter_out_expected[1423] <= 18'h0df04;
	 filter_out_expected[1424] <= 18'h2c6a4;
	 filter_out_expected[1425] <= 18'h1d4a3;
	 filter_out_expected[1426] <= 18'h31994;
	 filter_out_expected[1427] <= 18'h15e24;
	 filter_out_expected[1428] <= 18'h253bd;
	 filter_out_expected[1429] <= 18'h0f281;
	 filter_out_expected[1430] <= 18'h29252;
	 filter_out_expected[1431] <= 18'h195cb;
	 filter_out_expected[1432] <= 18'h2ff7e;
	 filter_out_expected[1433] <= 18'h169e0;
	 filter_out_expected[1434] <= 18'h26ee9;
	 filter_out_expected[1435] <= 18'h10f80;
	 filter_out_expected[1436] <= 18'h2ac19;
	 filter_out_expected[1437] <= 18'h19d01;
	 filter_out_expected[1438] <= 18'h2dfc3;
	 filter_out_expected[1439] <= 18'h12c40;
	 filter_out_expected[1440] <= 18'h2488a;
	 filter_out_expected[1441] <= 18'h134fd;
	 filter_out_expected[1442] <= 18'h30d13;
	 filter_out_expected[1443] <= 18'h1dd5c;
	 filter_out_expected[1444] <= 18'h2aeb1;
	 filter_out_expected[1445] <= 18'h0a7e9;
	 filter_out_expected[1446] <= 18'h1f5a6;
	 filter_out_expected[1447] <= 18'h179c1;
	 filter_out_expected[1448] <= 18'h3b44b;
	 filter_out_expected[1449] <= 18'h238a1;
	 filter_out_expected[1450] <= 18'h24c98;
	 filter_out_expected[1451] <= 18'h3e01a;
	 filter_out_expected[1452] <= 18'h19f3d;
	 filter_out_expected[1453] <= 18'h20320;
	 filter_out_expected[1454] <= 18'h09709;
	 filter_out_expected[1455] <= 18'h279d0;
	 filter_out_expected[1456] <= 18'h1936e;
	 filter_out_expected[1457] <= 18'h2ed07;
	 filter_out_expected[1458] <= 18'h18627;
	 filter_out_expected[1459] <= 18'h2f0db;
	 filter_out_expected[1460] <= 18'h189a0;
	 filter_out_expected[1461] <= 18'h2570b;
	 filter_out_expected[1462] <= 18'h072f3;
	 filter_out_expected[1463] <= 18'h2126b;
	 filter_out_expected[1464] <= 18'h1f685;
	 filter_out_expected[1465] <= 18'h038c1;
	 filter_out_expected[1466] <= 18'h22f0d;
	 filter_out_expected[1467] <= 18'h18d8e;
	 filter_out_expected[1468] <= 18'h31ac2;
	 filter_out_expected[1469] <= 18'h1c203;
	 filter_out_expected[1470] <= 18'h31947;
	 filter_out_expected[1471] <= 18'h17dc5;
	 filter_out_expected[1472] <= 18'h20d91;
	 filter_out_expected[1473] <= 18'h021e7;
	 filter_out_expected[1474] <= 18'h2164f;
	 filter_out_expected[1475] <= 18'h26760;
	 filter_out_expected[1476] <= 18'h0a982;
	 filter_out_expected[1477] <= 18'h210da;
	 filter_out_expected[1478] <= 18'h0e647;
	 filter_out_expected[1479] <= 18'h2a4d8;
	 filter_out_expected[1480] <= 18'h21de1;
	 filter_out_expected[1481] <= 18'h3f2db;
	 filter_out_expected[1482] <= 18'h1ced1;
	 filter_out_expected[1483] <= 18'h15ae5;
	 filter_out_expected[1484] <= 18'h33327;
	 filter_out_expected[1485] <= 18'h21ad3;
	 filter_out_expected[1486] <= 18'h37291;
	 filter_out_expected[1487] <= 18'h177ec;
	 filter_out_expected[1488] <= 18'h18f15;
	 filter_out_expected[1489] <= 18'h3a2cd;
	 filter_out_expected[1490] <= 18'h23a28;
	 filter_out_expected[1491] <= 18'h32815;
	 filter_out_expected[1492] <= 18'h12abe;
	 filter_out_expected[1493] <= 18'h199b4;
	 filter_out_expected[1494] <= 18'h3ea59;
	 filter_out_expected[1495] <= 18'h261b5;
	 filter_out_expected[1496] <= 18'h308a2;
	 filter_out_expected[1497] <= 18'h0f57e;
	 filter_out_expected[1498] <= 18'h18db4;
	 filter_out_expected[1499] <= 18'h00b73;
	 filter_out_expected[1500] <= 18'h28345;
	 filter_out_expected[1501] <= 18'h308f3;
	 filter_out_expected[1502] <= 18'h0db7a;
	 filter_out_expected[1503] <= 18'h17637;
	 filter_out_expected[1504] <= 18'h00b9b;
	 filter_out_expected[1505] <= 18'h29a79;
	 filter_out_expected[1506] <= 18'h3216f;
	 filter_out_expected[1507] <= 18'h0d9c2;
	 filter_out_expected[1508] <= 18'h156bc;
	 filter_out_expected[1509] <= 18'h3f0cb;
	 filter_out_expected[1510] <= 18'h2aa15;
	 filter_out_expected[1511] <= 18'h34e95;
	 filter_out_expected[1512] <= 18'h0e990;
	 filter_out_expected[1513] <= 18'h12cf4;
	 filter_out_expected[1514] <= 18'h3c125;
	 filter_out_expected[1515] <= 18'h2b9f3;
	 filter_out_expected[1516] <= 18'h38f22;
	 filter_out_expected[1517] <= 18'h100c7;
	 filter_out_expected[1518] <= 18'h0f36a;
	 filter_out_expected[1519] <= 18'h384a5;
	 filter_out_expected[1520] <= 18'h2d532;
	 filter_out_expected[1521] <= 18'h3e0cf;
	 filter_out_expected[1522] <= 18'h111cd;
	 filter_out_expected[1523] <= 18'h0a516;
	 filter_out_expected[1524] <= 18'h34774;
	 filter_out_expected[1525] <= 18'h3078e;
	 filter_out_expected[1526] <= 18'h03c5a;
	 filter_out_expected[1527] <= 18'h10c6d;
	 filter_out_expected[1528] <= 18'h04224;
	 filter_out_expected[1529] <= 18'h31b19;
	 filter_out_expected[1530] <= 18'h358b7;
	 filter_out_expected[1531] <= 18'h09232;
	 filter_out_expected[1532] <= 18'h0e1ac;
	 filter_out_expected[1533] <= 18'h3d524;
	 filter_out_expected[1534] <= 18'h3143b;
	 filter_out_expected[1535] <= 18'h3c597;
	 filter_out_expected[1536] <= 18'h0ca8c;
	 filter_out_expected[1537] <= 18'h08b73;
	 filter_out_expected[1538] <= 18'h375ca;
	 filter_out_expected[1539] <= 18'h342cf;
	 filter_out_expected[1540] <= 18'h03a46;
	 filter_out_expected[1541] <= 18'h0cc2d;
	 filter_out_expected[1542] <= 18'h01612;
	 filter_out_expected[1543] <= 18'h34490;
	 filter_out_expected[1544] <= 18'h3a579;
	 filter_out_expected[1545] <= 18'h0927d;
	 filter_out_expected[1546] <= 18'h08b22;
	 filter_out_expected[1547] <= 18'h3a4fb;
	 filter_out_expected[1548] <= 18'h35b7c;
	 filter_out_expected[1549] <= 18'h01ed5;
	 filter_out_expected[1550] <= 18'h0a752;
	 filter_out_expected[1551] <= 18'h019af;
	 filter_out_expected[1552] <= 18'h368e2;
	 filter_out_expected[1553] <= 18'h3b791;
	 filter_out_expected[1554] <= 18'h0792e;
	 filter_out_expected[1555] <= 18'h069e9;
	 filter_out_expected[1556] <= 18'h3acb2;
	 filter_out_expected[1557] <= 18'h38301;
	 filter_out_expected[1558] <= 18'h02aed;
	 filter_out_expected[1559] <= 18'h08280;
	 filter_out_expected[1560] <= 18'h3fb7f;
	 filter_out_expected[1561] <= 18'h38372;
	 filter_out_expected[1562] <= 18'h3e33c;
	 filter_out_expected[1563] <= 18'h06dff;
	 filter_out_expected[1564] <= 18'h036fa;
	 filter_out_expected[1565] <= 18'h3a622;
	 filter_out_expected[1566] <= 18'h3b69b;
	 filter_out_expected[1567] <= 18'h042fe;
	 filter_out_expected[1568] <= 18'h05435;
	 filter_out_expected[1569] <= 18'h3d43d;
	 filter_out_expected[1570] <= 18'h3a7bf;
	 filter_out_expected[1571] <= 18'h01600;
	 filter_out_expected[1572] <= 18'h056bf;
	 filter_out_expected[1573] <= 18'h3fd11;
	 filter_out_expected[1574] <= 18'h3aef2;
	 filter_out_expected[1575] <= 18'h3f343;
	 filter_out_expected[1576] <= 18'h0488a;
	 filter_out_expected[1577] <= 18'h018c4;
	 filter_out_expected[1578] <= 18'h3c196;
	 filter_out_expected[1579] <= 18'h3dec0;
	 filter_out_expected[1580] <= 18'h033ae;
	 filter_out_expected[1581] <= 18'h02680;
	 filter_out_expected[1582] <= 18'h3d6e0;
	 filter_out_expected[1583] <= 18'h3d709;
	 filter_out_expected[1584] <= 18'h01f50;
	 filter_out_expected[1585] <= 18'h0292b;
	 filter_out_expected[1586] <= 18'h3e968;
	 filter_out_expected[1587] <= 18'h3d864;
	 filter_out_expected[1588] <= 18'h00f26;
	 filter_out_expected[1589] <= 18'h024c3;
	 filter_out_expected[1590] <= 18'h3f6f6;
	 filter_out_expected[1591] <= 18'h3def6;
	 filter_out_expected[1592] <= 18'h00436;
	 filter_out_expected[1593] <= 18'h01cc6;
	 filter_out_expected[1594] <= 18'h3ff73;
	 filter_out_expected[1595] <= 18'h3e7c6;
	 filter_out_expected[1596] <= 18'h3fde9;
	 filter_out_expected[1597] <= 18'h01397;
	 filter_out_expected[1598] <= 18'h003e2;
	 filter_out_expected[1599] <= 18'h3f101;
	 filter_out_expected[1600] <= 18'h3fafd;
	 filter_out_expected[1601] <= 18'h00a8a;
	 filter_out_expected[1602] <= 18'h005a8;
	 filter_out_expected[1603] <= 18'h3f9bc;
	 filter_out_expected[1604] <= 18'h3fa04;
	 filter_out_expected[1605] <= 18'h00234;
	 filter_out_expected[1606] <= 18'h00628;
	 filter_out_expected[1607] <= 18'h001a4;
	 filter_out_expected[1608] <= 18'h3f9af;
	 filter_out_expected[1609] <= 18'h3fabd;
	 filter_out_expected[1610] <= 18'h00699;
	 filter_out_expected[1611] <= 18'h008a7;
	 filter_out_expected[1612] <= 18'h3f8e4;
	 filter_out_expected[1613] <= 18'h3f437;
	 filter_out_expected[1614] <= 18'h007f9;
	 filter_out_expected[1615] <= 18'h00ea2;
	 filter_out_expected[1616] <= 18'h3f6bd;
	 filter_out_expected[1617] <= 18'h3eedb;
	 filter_out_expected[1618] <= 18'h00b0c;
	 filter_out_expected[1619] <= 18'h0133a;
	 filter_out_expected[1620] <= 18'h3f2a1;
	 filter_out_expected[1621] <= 18'h3eb37;
	 filter_out_expected[1622] <= 18'h0103e;
	 filter_out_expected[1623] <= 18'h015b0;
	 filter_out_expected[1624] <= 18'h3ec5d;
	 filter_out_expected[1625] <= 18'h3ea37;
	 filter_out_expected[1626] <= 18'h01778;
	 filter_out_expected[1627] <= 18'h014ec;
	 filter_out_expected[1628] <= 18'h3e465;
	 filter_out_expected[1629] <= 18'h3ed10;
	 filter_out_expected[1630] <= 18'h01fd9;
	 filter_out_expected[1631] <= 18'h00fb3;
	 filter_out_expected[1632] <= 18'h3dc15;
	 filter_out_expected[1633] <= 18'h3f4e3;
	 filter_out_expected[1634] <= 18'h0277b;
	 filter_out_expected[1635] <= 18'h00529;
	 filter_out_expected[1636] <= 18'h3d5de;
	 filter_out_expected[1637] <= 18'h00214;
	 filter_out_expected[1638] <= 18'h02b6f;
	 filter_out_expected[1639] <= 18'h3f59a;
	 filter_out_expected[1640] <= 18'h3d50d;
	 filter_out_expected[1641] <= 18'h0136f;
	 filter_out_expected[1642] <= 18'h02844;
	 filter_out_expected[1643] <= 18'h3e358;
	 filter_out_expected[1644] <= 18'h3dceb;
	 filter_out_expected[1645] <= 18'h02562;
	 filter_out_expected[1646] <= 18'h01b42;
	 filter_out_expected[1647] <= 18'h3d337;
	 filter_out_expected[1648] <= 18'h3ef1d;
	 filter_out_expected[1649] <= 18'h031f6;
	 filter_out_expected[1650] <= 18'h0045e;
	 filter_out_expected[1651] <= 18'h3cbfa;
	 filter_out_expected[1652] <= 18'h00990;
	 filter_out_expected[1653] <= 18'h03238;
	 filter_out_expected[1654] <= 18'h3e82e;
	 filter_out_expected[1655] <= 18'h3d3ef;
	 filter_out_expected[1656] <= 18'h02509;
	 filter_out_expected[1657] <= 18'h02180;
	 filter_out_expected[1658] <= 18'h3d05d;
	 filter_out_expected[1659] <= 18'h3ecfd;
	 filter_out_expected[1660] <= 18'h03612;
	 filter_out_expected[1661] <= 18'h001b7;
	 filter_out_expected[1662] <= 18'h3c900;
	 filter_out_expected[1663] <= 18'h010ab;
	 filter_out_expected[1664] <= 18'h0319a;
	 filter_out_expected[1665] <= 18'h3de18;
	 filter_out_expected[1666] <= 18'h3da2a;
	 filter_out_expected[1667] <= 18'h02f88;
	 filter_out_expected[1668] <= 18'h0149e;
	 filter_out_expected[1669] <= 18'h3c8ce;
	 filter_out_expected[1670] <= 18'h00018;
	 filter_out_expected[1671] <= 18'h03720;
	 filter_out_expected[1672] <= 18'h3ea94;
	 filter_out_expected[1673] <= 18'h3d166;
	 filter_out_expected[1674] <= 18'h027f0;
	 filter_out_expected[1675] <= 18'h01e4d;
	 filter_out_expected[1676] <= 18'h3cbce;
	 filter_out_expected[1677] <= 18'h3f78c;
	 filter_out_expected[1678] <= 18'h03778;
	 filter_out_expected[1679] <= 18'h3f0b2;
	 filter_out_expected[1680] <= 18'h3cf89;
	 filter_out_expected[1681] <= 18'h02474;
	 filter_out_expected[1682] <= 18'h01fde;
	 filter_out_expected[1683] <= 18'h3cd87;
	 filter_out_expected[1684] <= 18'h3f773;
	 filter_out_expected[1685] <= 18'h035ea;
	 filter_out_expected[1686] <= 18'h3ef45;
	 filter_out_expected[1687] <= 18'h3d29d;
	 filter_out_expected[1688] <= 18'h02641;
	 filter_out_expected[1689] <= 18'h01a4a;
	 filter_out_expected[1690] <= 18'h3cd5f;
	 filter_out_expected[1691] <= 18'h3ff2a;
	 filter_out_expected[1692] <= 18'h03250;
	 filter_out_expected[1693] <= 18'h3e753;
	 filter_out_expected[1694] <= 18'h3db21;
	 filter_out_expected[1695] <= 18'h02b61;
	 filter_out_expected[1696] <= 18'h00d88;
	 filter_out_expected[1697] <= 18'h3ce39;
	 filter_out_expected[1698] <= 18'h00d55;
	 filter_out_expected[1699] <= 18'h029a1;
	 filter_out_expected[1700] <= 18'h3dc32;
	 filter_out_expected[1701] <= 18'h3eaf4;
	 filter_out_expected[1702] <= 18'h02ec9;
	 filter_out_expected[1703] <= 18'h3fa48;
	 filter_out_expected[1704] <= 18'h3d57f;
	 filter_out_expected[1705] <= 18'h01df9;
	 filter_out_expected[1706] <= 18'h01829;
	 filter_out_expected[1707] <= 18'h3d4a1;
	 filter_out_expected[1708] <= 18'h00206;
	 filter_out_expected[1709] <= 18'h02912;
	 filter_out_expected[1710] <= 18'h3e559;
	 filter_out_expected[1711] <= 18'h3e82f;
	 filter_out_expected[1712] <= 18'h0287e;
	 filter_out_expected[1713] <= 18'h3fe29;
	 filter_out_expected[1714] <= 18'h3d9d1;
	 filter_out_expected[1715] <= 18'h019c2;
	 filter_out_expected[1716] <= 18'h014b7;
	 filter_out_expected[1717] <= 18'h3d9cf;
	 filter_out_expected[1718] <= 18'h00488;
	 filter_out_expected[1719] <= 18'h02203;
	 filter_out_expected[1720] <= 18'h3e55c;
	 filter_out_expected[1721] <= 18'h3f0b9;
	 filter_out_expected[1722] <= 18'h023e0;
	 filter_out_expected[1723] <= 18'h3f6b1;
	 filter_out_expected[1724] <= 18'h3e3ba;
	 filter_out_expected[1725] <= 18'h01c36;
	 filter_out_expected[1726] <= 18'h007d9;
	 filter_out_expected[1727] <= 18'h3df78;
	 filter_out_expected[1728] <= 18'h00f1c;
	 filter_out_expected[1729] <= 18'h0149a;
	 filter_out_expected[1730] <= 18'h3e2f9;
	 filter_out_expected[1731] <= 18'h000ef;
	 filter_out_expected[1732] <= 18'h01b16;
	 filter_out_expected[1733] <= 18'h3eb92;
	 filter_out_expected[1734] <= 18'h3f501;
	 filter_out_expected[1735] <= 18'h01b82;
	 filter_out_expected[1736] <= 18'h3f636;
	 filter_out_expected[1737] <= 18'h3ed1b;
	 filter_out_expected[1738] <= 18'h01762;
	 filter_out_expected[1739] <= 18'h0005b;
	 filter_out_expected[1740] <= 18'h3e998;
	 filter_out_expected[1741] <= 18'h010b2;
	 filter_out_expected[1742] <= 18'h00861;
	 filter_out_expected[1743] <= 18'h3e9d2;
	 filter_out_expected[1744] <= 18'h00949;
	 filter_out_expected[1745] <= 18'h00d9b;
	 filter_out_expected[1746] <= 18'h3eca5;
	 filter_out_expected[1747] <= 18'h00283;
	 filter_out_expected[1748] <= 18'h01017;
	 filter_out_expected[1749] <= 18'h3f0dc;
	 filter_out_expected[1750] <= 18'h3fd27;
	 filter_out_expected[1751] <= 18'h01056;
	 filter_out_expected[1752] <= 18'h3f570;
	 filter_out_expected[1753] <= 18'h3f97f;
	 filter_out_expected[1754] <= 18'h00f05;
	 filter_out_expected[1755] <= 18'h3f9ab;
	 filter_out_expected[1756] <= 18'h3f778;
	 filter_out_expected[1757] <= 18'h00cd0;
	 filter_out_expected[1758] <= 18'h3fd23;
	 filter_out_expected[1759] <= 18'h3f6cd;
	 filter_out_expected[1760] <= 18'h00a40;
	 filter_out_expected[1761] <= 18'h3ffaf;
	 filter_out_expected[1762] <= 18'h3f722;
	 filter_out_expected[1763] <= 18'h007b7;
	 filter_out_expected[1764] <= 18'h00154;
	 filter_out_expected[1765] <= 18'h3f824;
	 filter_out_expected[1766] <= 18'h00571;
	 filter_out_expected[1767] <= 18'h00233;
	 filter_out_expected[1768] <= 18'h3f98a;
	 filter_out_expected[1769] <= 18'h00385;
	 filter_out_expected[1770] <= 18'h00275;
	 filter_out_expected[1771] <= 18'h3fb20;
	 filter_out_expected[1772] <= 18'h001f5;
	 filter_out_expected[1773] <= 18'h00247;
	 filter_out_expected[1774] <= 18'h3fcc2;
	 filter_out_expected[1775] <= 18'h000b4;
	 filter_out_expected[1776] <= 18'h001d4;
	 filter_out_expected[1777] <= 18'h3fe5d;
	 filter_out_expected[1778] <= 18'h3ffac;
	 filter_out_expected[1779] <= 18'h00140;
	 filter_out_expected[1780] <= 18'h3ffe5;
	 filter_out_expected[1781] <= 18'h3fec2;
	 filter_out_expected[1782] <= 18'h000ab;
	 filter_out_expected[1783] <= 18'h00155;
	 filter_out_expected[1784] <= 18'h3fde0;
	 filter_out_expected[1785] <= 18'h00032;
	 filter_out_expected[1786] <= 18'h002aa;
	 filter_out_expected[1787] <= 18'h3fcef;
	 filter_out_expected[1788] <= 18'h3fff1;
	 filter_out_expected[1789] <= 18'h003d8;
	 filter_out_expected[1790] <= 18'h3fbdf;
	 filter_out_expected[1791] <= 18'h3fffd;
	 filter_out_expected[1792] <= 18'h004d2;
	 filter_out_expected[1793] <= 18'h3faac;
	 filter_out_expected[1794] <= 18'h0006f;
	 filter_out_expected[1795] <= 18'h00583;
	 filter_out_expected[1796] <= 18'h3f95a;
	 filter_out_expected[1797] <= 18'h0015a;
	 filter_out_expected[1798] <= 18'h005ca;
	 filter_out_expected[1799] <= 18'h3f7ff;
	 filter_out_expected[1800] <= 18'h002c5;
	 filter_out_expected[1801] <= 18'h00582;
	 filter_out_expected[1802] <= 18'h3f6c1;
	 filter_out_expected[1803] <= 18'h004a9;
	 filter_out_expected[1804] <= 18'h00485;
	 filter_out_expected[1805] <= 18'h3f5da;
	 filter_out_expected[1806] <= 18'h006ea;
	 filter_out_expected[1807] <= 18'h002b6;
	 filter_out_expected[1808] <= 18'h3f594;
	 filter_out_expected[1809] <= 18'h00949;
	 filter_out_expected[1810] <= 18'h0000d;
	 filter_out_expected[1811] <= 18'h3f63f;
	 filter_out_expected[1812] <= 18'h00b6c;
	 filter_out_expected[1813] <= 18'h3fca9;
	 filter_out_expected[1814] <= 18'h3f81e;
	 filter_out_expected[1815] <= 18'h00cd2;
	 filter_out_expected[1816] <= 18'h3f8db;
	 filter_out_expected[1817] <= 18'h3fb55;
	 filter_out_expected[1818] <= 18'h00cf5;
	 filter_out_expected[1819] <= 18'h3f532;
	 filter_out_expected[1820] <= 18'h3ffc5;
	 filter_out_expected[1821] <= 18'h00b58;
	 filter_out_expected[1822] <= 18'h3f270;
	 filter_out_expected[1823] <= 18'h004f9;
	 filter_out_expected[1824] <= 18'h007bd;
	 filter_out_expected[1825] <= 18'h3f16d;
	 filter_out_expected[1826] <= 18'h00a18;
	 filter_out_expected[1827] <= 18'h0024f;
	 filter_out_expected[1828] <= 18'h3f2e5;
	 filter_out_expected[1829] <= 18'h00dfb;
	 filter_out_expected[1830] <= 18'h3fbcc;
	 filter_out_expected[1831] <= 18'h3f722;
	 filter_out_expected[1832] <= 18'h00f63;
	 filter_out_expected[1833] <= 18'h3f587;
	 filter_out_expected[1834] <= 18'h3fdc0;
	 filter_out_expected[1835] <= 18'h00d66;
	 filter_out_expected[1836] <= 18'h3f133;
	 filter_out_expected[1837] <= 18'h00575;
	 filter_out_expected[1838] <= 18'h007db;
	 filter_out_expected[1839] <= 18'h3f06d;
	 filter_out_expected[1840] <= 18'h00c38;
	 filter_out_expected[1841] <= 18'h3ffc5;
	 filter_out_expected[1842] <= 18'h3f414;
	 filter_out_expected[1843] <= 18'h00fbf;
	 filter_out_expected[1844] <= 18'h3f755;
	 filter_out_expected[1845] <= 18'h3fba9;
	 filter_out_expected[1846] <= 18'h00e58;
	 filter_out_expected[1847] <= 18'h3f16b;
	 filter_out_expected[1848] <= 18'h00503;
	 filter_out_expected[1849] <= 18'h007d8;
	 filter_out_expected[1850] <= 18'h3f098;
	 filter_out_expected[1851] <= 18'h00cc4;
	 filter_out_expected[1852] <= 18'h3fe32;
	 filter_out_expected[1853] <= 18'h3f5c8;
	 filter_out_expected[1854] <= 18'h00f88;
	 filter_out_expected[1855] <= 18'h3f525;
	 filter_out_expected[1856] <= 18'h3ff58;
	 filter_out_expected[1857] <= 18'h00b9b;
	 filter_out_expected[1858] <= 18'h3f0db;
	 filter_out_expected[1859] <= 18'h0093a;
	 filter_out_expected[1860] <= 18'h0024a;
	 filter_out_expected[1861] <= 18'h3f3ca;
	 filter_out_expected[1862] <= 18'h00e8e;
	 filter_out_expected[1863] <= 18'h3f7ec;
	 filter_out_expected[1864] <= 18'h3fce5;
	 filter_out_expected[1865] <= 18'h00c3a;
	 filter_out_expected[1866] <= 18'h3f209;
	 filter_out_expected[1867] <= 18'h0077e;
	 filter_out_expected[1868] <= 18'h0032e;
	 filter_out_expected[1869] <= 18'h3f439;
	 filter_out_expected[1870] <= 18'h00d72;
	 filter_out_expected[1871] <= 18'h3f88f;
	 filter_out_expected[1872] <= 18'h3fd68;
	 filter_out_expected[1873] <= 18'h00aea;
	 filter_out_expected[1874] <= 18'h3f309;
	 filter_out_expected[1875] <= 18'h007d5;
	 filter_out_expected[1876] <= 18'h0016c;
	 filter_out_expected[1877] <= 18'h3f65f;
	 filter_out_expected[1878] <= 18'h00c6a;
	 filter_out_expected[1879] <= 18'h3f780;
	 filter_out_expected[1880] <= 18'h0003b;
	 filter_out_expected[1881] <= 18'h007e2;
	 filter_out_expected[1882] <= 18'h3f463;
	 filter_out_expected[1883] <= 18'h0093a;
	 filter_out_expected[1884] <= 18'h3fdca;
	 filter_out_expected[1885] <= 18'h3fa58;
	 filter_out_expected[1886] <= 18'h00a5f;
	 filter_out_expected[1887] <= 18'h3f647;
	 filter_out_expected[1888] <= 18'h0044c;
	 filter_out_expected[1889] <= 18'h00302;
	 filter_out_expected[1890] <= 18'h3f77a;
	 filter_out_expected[1891] <= 18'h009ae;
	 filter_out_expected[1892] <= 18'h3f9d8;
	 filter_out_expected[1893] <= 18'h3ffe3;
	 filter_out_expected[1894] <= 18'h00605;
	 filter_out_expected[1895] <= 18'h3f72e;
	 filter_out_expected[1896] <= 18'h00766;
	 filter_out_expected[1897] <= 18'h3fd55;
	 filter_out_expected[1898] <= 18'h3fcff;
	 filter_out_expected[1899] <= 18'h00701;
	 filter_out_expected[1900] <= 18'h3f85c;
	 filter_out_expected[1901] <= 18'h004dd;
	 filter_out_expected[1902] <= 18'h3ffdd;
	 filter_out_expected[1903] <= 18'h3fba8;
	 filter_out_expected[1904] <= 18'h006a6;
	 filter_out_expected[1905] <= 18'h3fa0a;
	 filter_out_expected[1906] <= 18'h002cf;
	 filter_out_expected[1907] <= 18'h00149;
	 filter_out_expected[1908] <= 18'h3fb7b;
	 filter_out_expected[1909] <= 18'h005a4;
	 filter_out_expected[1910] <= 18'h3fba1;
	 filter_out_expected[1911] <= 18'h00173;
	 filter_out_expected[1912] <= 18'h001c7;
	 filter_out_expected[1913] <= 18'h3fc00;
	 filter_out_expected[1914] <= 18'h0046e;
	 filter_out_expected[1915] <= 18'h3fce8;
	 filter_out_expected[1916] <= 18'h000b8;
	 filter_out_expected[1917] <= 18'h001aa;
	 filter_out_expected[1918] <= 18'h3fce1;
	 filter_out_expected[1919] <= 18'h00339;
	 filter_out_expected[1920] <= 18'h3fde3;
	 filter_out_expected[1921] <= 18'h00062;
	 filter_out_expected[1922] <= 18'h00138;
	 filter_out_expected[1923] <= 18'h3fde4;
	 filter_out_expected[1924] <= 18'h00212;
	 filter_out_expected[1925] <= 18'h3feb6;
	 filter_out_expected[1926] <= 18'h00034;
	 filter_out_expected[1927] <= 18'h000b4;
	 filter_out_expected[1928] <= 18'h3fee4;
	 filter_out_expected[1929] <= 18'h000f7;
	 filter_out_expected[1930] <= 18'h3ff89;
	 filter_out_expected[1931] <= 18'h3fff0;
	 filter_out_expected[1932] <= 18'h0005a;
	 filter_out_expected[1933] <= 18'h3ffb9;
	 filter_out_expected[1934] <= 18'h3ffee;
	 filter_out_expected[1935] <= 18'h00073;
	 filter_out_expected[1936] <= 18'h3ff64;
	 filter_out_expected[1937] <= 18'h00063;
	 filter_out_expected[1938] <= 18'h00030;
	 filter_out_expected[1939] <= 18'h3ff1c;
	 filter_out_expected[1940] <= 18'h0016d;
	 filter_out_expected[1941] <= 18'h3fe7f;
	 filter_out_expected[1942] <= 18'h000fd;
	 filter_out_expected[1943] <= 18'h00002;
	 filter_out_expected[1944] <= 18'h3fecb;
	 filter_out_expected[1945] <= 18'h00231;
	 filter_out_expected[1946] <= 18'h3fd6b;
	 filter_out_expected[1947] <= 18'h0022b;
	 filter_out_expected[1948] <= 18'h3ff01;
	 filter_out_expected[1949] <= 18'h3ff5c;
	 filter_out_expected[1950] <= 18'h00243;
	 filter_out_expected[1951] <= 18'h3fca4;
	 filter_out_expected[1952] <= 18'h0038f;
	 filter_out_expected[1953] <= 18'h3fd47;
	 filter_out_expected[1954] <= 18'h00108;
	 filter_out_expected[1955] <= 18'h00118;
	 filter_out_expected[1956] <= 18'h3fcef;
	 filter_out_expected[1957] <= 18'h00454;
	 filter_out_expected[1958] <= 18'h3fb82;
	 filter_out_expected[1959] <= 18'h00377;
	 filter_out_expected[1960] <= 18'h3fe8c;
	 filter_out_expected[1961] <= 18'h3fef5;
	 filter_out_expected[1962] <= 18'h00366;
	 filter_out_expected[1963] <= 18'h3fafd;
	 filter_out_expected[1964] <= 18'h00571;
	 filter_out_expected[1965] <= 18'h3fb74;
	 filter_out_expected[1966] <= 18'h00284;
	 filter_out_expected[1967] <= 18'h00035;
	 filter_out_expected[1968] <= 18'h3fd07;
	 filter_out_expected[1969] <= 18'h00524;
	 filter_out_expected[1970] <= 18'h3f9cd;
	 filter_out_expected[1971] <= 18'h005e0;
	 filter_out_expected[1972] <= 18'h3fbc5;
	 filter_out_expected[1973] <= 18'h0019b;
	 filter_out_expected[1974] <= 18'h00170;
	 filter_out_expected[1975] <= 18'h3fbc3;
	 filter_out_expected[1976] <= 18'h00635;
	 filter_out_expected[1977] <= 18'h3f915;
	 filter_out_expected[1978] <= 18'h00637;
	 filter_out_expected[1979] <= 18'h3fbc3;
	 filter_out_expected[1980] <= 18'h00161;
	 filter_out_expected[1981] <= 18'h001cd;
	 filter_out_expected[1982] <= 18'h3fb55;
	 filter_out_expected[1983] <= 18'h006ad;
	 filter_out_expected[1984] <= 18'h3f88d;
	 filter_out_expected[1985] <= 18'h006d4;
	 filter_out_expected[1986] <= 18'h3fb0c;
	 filter_out_expected[1987] <= 18'h00229;
	 filter_out_expected[1988] <= 18'h0010a;
	 filter_out_expected[1989] <= 18'h3fbee;
	 filter_out_expected[1990] <= 18'h0066a;
	 filter_out_expected[1991] <= 18'h3f854;
	 filter_out_expected[1992] <= 18'h007a2;
	 filter_out_expected[1993] <= 18'h3f9ab;
	 filter_out_expected[1994] <= 18'h003fe;
	 filter_out_expected[1995] <= 18'h3fefe;
	 filter_out_expected[1996] <= 18'h3fdde;
	 filter_out_expected[1997] <= 18'h004ef;
	 filter_out_expected[1998] <= 18'h3f908;
	 filter_out_expected[1999] <= 18'h007f1;
	 filter_out_expected[2000] <= 18'h3f846;
	 filter_out_expected[2001] <= 18'h00661;
	 filter_out_expected[2002] <= 18'h3fbe2;
	 filter_out_expected[2003] <= 18'h00149;
	 filter_out_expected[2004] <= 18'h001b4;
	 filter_out_expected[2005] <= 18'h3fb91;
	 filter_out_expected[2006] <= 18'h00689;
	 filter_out_expected[2007] <= 18'h3f841;
	 filter_out_expected[2008] <= 18'h007ee;
	 filter_out_expected[2009] <= 18'h3f8ea;
	 filter_out_expected[2010] <= 18'h0055c;
	 filter_out_expected[2011] <= 18'h3fd03;
	 filter_out_expected[2012] <= 18'h00048;
	 filter_out_expected[2013] <= 18'h0026a;
	 filter_out_expected[2014] <= 18'h3fb37;
	 filter_out_expected[2015] <= 18'h0068f;
	 filter_out_expected[2016] <= 18'h3f872;
	 filter_out_expected[2017] <= 18'h007ae;
	 filter_out_expected[2018] <= 18'h3f909;
	 filter_out_expected[2019] <= 18'h00581;
	 filter_out_expected[2020] <= 18'h3fc82;
	 filter_out_expected[2021] <= 18'h00129;
	 filter_out_expected[2022] <= 18'h0013e;
	 filter_out_expected[2023] <= 18'h3fc89;
	 filter_out_expected[2024] <= 18'h0054a;
	 filter_out_expected[2025] <= 18'h3f970;
	 filter_out_expected[2026] <= 18'h0072d;
	 filter_out_expected[2027] <= 18'h3f8e4;
	 filter_out_expected[2028] <= 18'h00666;
	 filter_out_expected[2029] <= 18'h3fadf;
	 filter_out_expected[2030] <= 18'h00373;
	 filter_out_expected[2031] <= 18'h3fe7a;
	 filter_out_expected[2032] <= 18'h3ff86;
	 filter_out_expected[2033] <= 18'h0025f;
	 filter_out_expected[2034] <= 18'h3fbfc;
	 filter_out_expected[2035] <= 18'h0054a;
	 filter_out_expected[2036] <= 18'h3f9e4;
	 filter_out_expected[2037] <= 18'h00671;
	 filter_out_expected[2038] <= 18'h3f9b9;
	 filter_out_expected[2039] <= 18'h005ab;
	 filter_out_expected[2040] <= 18'h3fb52;
	 filter_out_expected[2041] <= 18'h00366;
	 filter_out_expected[2042] <= 18'h3fe0f;
	 filter_out_expected[2043] <= 18'h00068;
	 filter_out_expected[2044] <= 18'h00116;
	 filter_out_expected[2045] <= 18'h3fd8c;
	 filter_out_expected[2046] <= 18'h0039c;
	 filter_out_expected[2047] <= 18'h3fb82;
	 filter_out_expected[2048] <= 18'h00514;
	 filter_out_expected[2049] <= 18'h3faa9;
	 filter_out_expected[2050] <= 18'h0054a;
	 filter_out_expected[2051] <= 18'h3fb0d;
	 filter_out_expected[2052] <= 18'h0045c;
	 filter_out_expected[2053] <= 18'h3fc6d;
	 filter_out_expected[2054] <= 18'h002a4;
	 filter_out_expected[2055] <= 18'h3fe60;
	 filter_out_expected[2056] <= 18'h00096;
	 filter_out_expected[2057] <= 18'h0006e;
	 filter_out_expected[2058] <= 18'h3fea2;
	 filter_out_expected[2059] <= 18'h00231;
	 filter_out_expected[2060] <= 18'h3fd21;
	 filter_out_expected[2061] <= 18'h00364;
	 filter_out_expected[2062] <= 18'h3fc42;
	 filter_out_expected[2063] <= 18'h003eb;
	 filter_out_expected[2064] <= 18'h3fc12;
	 filter_out_expected[2065] <= 18'h003cb;
	 filter_out_expected[2066] <= 18'h3fc7a;
	 filter_out_expected[2067] <= 18'h00324;
	 filter_out_expected[2068] <= 18'h3fd53;
	 filter_out_expected[2069] <= 18'h00227;
	 filter_out_expected[2070] <= 18'h3fe68;
	 filter_out_expected[2071] <= 18'h00106;
	 filter_out_expected[2072] <= 18'h3ff8a;
	 filter_out_expected[2073] <= 18'h3ffed;
	 filter_out_expected[2074] <= 18'h00091;
	 filter_out_expected[2075] <= 18'h3feff;
	 filter_out_expected[2076] <= 18'h00161;
	 filter_out_expected[2077] <= 18'h3fe51;
	 filter_out_expected[2078] <= 18'h001ec;
	 filter_out_expected[2079] <= 18'h3fde8;
	 filter_out_expected[2080] <= 18'h00232;
	 filter_out_expected[2081] <= 18'h3fdc4;
	 filter_out_expected[2082] <= 18'h00238;
	 filter_out_expected[2083] <= 18'h3fdd9;
	 filter_out_expected[2084] <= 18'h0020c;
	 filter_out_expected[2085] <= 18'h3fe19;
	 filter_out_expected[2086] <= 18'h001bc;
	 filter_out_expected[2087] <= 18'h3fe73;
	 filter_out_expected[2088] <= 18'h00158;
	 filter_out_expected[2089] <= 18'h3fedc;
	 filter_out_expected[2090] <= 18'h000ef;
	 filter_out_expected[2091] <= 18'h3ff46;
	 filter_out_expected[2092] <= 18'h00089;
	 filter_out_expected[2093] <= 18'h3ffa7;
	 filter_out_expected[2094] <= 18'h0002e;
	 filter_out_expected[2095] <= 18'h3fff9;
	 filter_out_expected[2096] <= 18'h3ffe4;
	 filter_out_expected[2097] <= 18'h0003b;
	 filter_out_expected[2098] <= 18'h3ffab;
	 filter_out_expected[2099] <= 18'h0006b;
	 filter_out_expected[2100] <= 18'h3ff84;
	 filter_out_expected[2101] <= 18'h0008a;
	 filter_out_expected[2102] <= 18'h3ff6d;
	 filter_out_expected[2103] <= 18'h0227d;
	 filter_out_expected[2104] <= 18'h035f2;
	 filter_out_expected[2105] <= 18'h02103;
	 filter_out_expected[2106] <= 18'h3dceb;
	 filter_out_expected[2107] <= 18'h3a8aa;
	 filter_out_expected[2108] <= 18'h3a804;
	 filter_out_expected[2109] <= 18'h3e123;
	 filter_out_expected[2110] <= 18'h02117;
	 filter_out_expected[2111] <= 18'h03749;
	 filter_out_expected[2112] <= 18'h01fbe;
	 filter_out_expected[2113] <= 18'h00000;
	 filter_out_expected[2114] <= 18'h01ea9;
	 filter_out_expected[2115] <= 18'h07d70;
	 filter_out_expected[2116] <= 18'h0b0ce;
	 filter_out_expected[2117] <= 18'h049fb;
	 filter_out_expected[2118] <= 18'h36e15;
	 filter_out_expected[2119] <= 18'h2c56c;
	 filter_out_expected[2120] <= 18'h2dd96;
	 filter_out_expected[2121] <= 18'h3c779;
	 filter_out_expected[2122] <= 18'h0bd30;
	 filter_out_expected[2123] <= 18'h0ae62;
	 filter_out_expected[2124] <= 18'h3b640;
	 filter_out_expected[2125] <= 18'h2df9a;
	 filter_out_expected[2126] <= 18'h32d0d;
	 filter_out_expected[2127] <= 18'h05958;
	 filter_out_expected[2128] <= 18'h16742;
	 filter_out_expected[2129] <= 18'h186a8;
	 filter_out_expected[2130] <= 18'h0cd7a;
	 filter_out_expected[2131] <= 18'h01da5;
	 filter_out_expected[2132] <= 18'h3f8d3;
	 filter_out_expected[2133] <= 18'h01570;
	 filter_out_expected[2134] <= 18'h3c5c3;
	 filter_out_expected[2135] <= 18'h2e9d3;
	 filter_out_expected[2136] <= 18'h25bb1;
	 filter_out_expected[2137] <= 18'h30117;
	 filter_out_expected[2138] <= 18'h09035;
	 filter_out_expected[2139] <= 18'h1a1c5;
	 filter_out_expected[2140] <= 18'h10e59;
	 filter_out_expected[2141] <= 18'h39041;
	 filter_out_expected[2142] <= 18'h29f56;
	 filter_out_expected[2143] <= 18'h31fdc;
	 filter_out_expected[2144] <= 18'h08d5d;
	 filter_out_expected[2145] <= 18'h13dea;
	 filter_out_expected[2146] <= 18'h07bd9;
	 filter_out_expected[2147] <= 18'h34184;
	 filter_out_expected[2148] <= 18'h2b013;
	 filter_out_expected[2149] <= 18'h31827;
	 filter_out_expected[2150] <= 18'h049cc;
	 filter_out_expected[2151] <= 18'h188fe;
	 filter_out_expected[2152] <= 18'h24356;
	 filter_out_expected[2153] <= 18'h1fc6d;
	 filter_out_expected[2154] <= 18'h0d6d6;
	 filter_out_expected[2155] <= 18'h357b2;
	 filter_out_expected[2156] <= 18'h1d0b0;
	 filter_out_expected[2157] <= 18'h12cdf;
	 filter_out_expected[2158] <= 18'h1ee9e;
	 filter_out_expected[2159] <= 18'h364f6;
	 filter_out_expected[2160] <= 18'h07883;
	 filter_out_expected[2161] <= 18'h0b999;
	 filter_out_expected[2162] <= 18'h05b0c;
	 filter_out_expected[2163] <= 18'h3f875;
	 filter_out_expected[2164] <= 18'h05b1b;
	 filter_out_expected[2165] <= 18'h14c3e;
	 filter_out_expected[2166] <= 18'h1cde5;
	 filter_out_expected[2167] <= 18'h16a87;
	 filter_out_expected[2168] <= 18'h07a16;
	 filter_out_expected[2169] <= 18'h3793d;
	 filter_out_expected[2170] <= 18'h2bdd5;
	 filter_out_expected[2171] <= 18'h2a191;
	 filter_out_expected[2172] <= 18'h31798;
	 filter_out_expected[2173] <= 18'h3a244;
	 filter_out_expected[2174] <= 18'h3fbad;
	 filter_out_expected[2175] <= 18'h03c42;
	 filter_out_expected[2176] <= 18'h0689c;
	 filter_out_expected[2177] <= 18'h0afd3;
	 filter_out_expected[2178] <= 18'h0e624;
	 filter_out_expected[2179] <= 18'h0520a;
	 filter_out_expected[2180] <= 18'h34600;
	 filter_out_expected[2181] <= 18'h2aa28;
	 filter_out_expected[2182] <= 18'h2fc62;
	 filter_out_expected[2183] <= 18'h3eb06;
	 filter_out_expected[2184] <= 18'h0c36d;
	 filter_out_expected[2185] <= 18'h11ad0;
	 filter_out_expected[2186] <= 18'h0f667;
	 filter_out_expected[2187] <= 18'h0d289;
	 filter_out_expected[2188] <= 18'h0cb7f;
	 filter_out_expected[2189] <= 18'h04a67;
	 filter_out_expected[2190] <= 18'h2f8e1;
	 filter_out_expected[2191] <= 18'h1cf73;
	 filter_out_expected[2192] <= 18'h20622;
	 filter_out_expected[2193] <= 18'h39192;
	 filter_out_expected[2194] <= 18'h0f3ee;
	 filter_out_expected[2195] <= 18'h0f70b;
	 filter_out_expected[2196] <= 18'h04083;
	 filter_out_expected[2197] <= 18'h0186d;
	 filter_out_expected[2198] <= 18'h0a888;
	 filter_out_expected[2199] <= 18'h0f588;
	 filter_out_expected[2200] <= 18'h05a89;
	 filter_out_expected[2201] <= 18'h37f5d;
	 filter_out_expected[2202] <= 18'h344c0;
	 filter_out_expected[2203] <= 18'h3cd16;
	 filter_out_expected[2204] <= 18'h03124;
	 filter_out_expected[2205] <= 18'h3ebf8;
	 filter_out_expected[2206] <= 18'h3bf2e;
	 filter_out_expected[2207] <= 18'h0127c;
	 filter_out_expected[2208] <= 18'h039ca;
	 filter_out_expected[2209] <= 18'h383e5;
	 filter_out_expected[2210] <= 18'h2ce56;
	 filter_out_expected[2211] <= 18'h37540;
	 filter_out_expected[2212] <= 18'h146c7;
	 filter_out_expected[2213] <= 18'h2748f;
	 filter_out_expected[2214] <= 18'h1c356;
	 filter_out_expected[2215] <= 18'h3a308;
	 filter_out_expected[2216] <= 18'h1dc1a;
	 filter_out_expected[2217] <= 18'h2191e;
	 filter_out_expected[2218] <= 18'h3b305;
	 filter_out_expected[2219] <= 18'h0c294;
	 filter_out_expected[2220] <= 18'h06cda;
	 filter_out_expected[2221] <= 18'h3ae99;
	 filter_out_expected[2222] <= 18'h3a715;
	 filter_out_expected[2223] <= 18'h05e33;
	 filter_out_expected[2224] <= 18'h0eead;
	 filter_out_expected[2225] <= 18'h0648c;
	 filter_out_expected[2226] <= 18'h2f643;
	 filter_out_expected[2227] <= 18'h24b12;
	 filter_out_expected[2228] <= 18'h36ad8;
	 filter_out_expected[2229] <= 18'h14314;
	 filter_out_expected[2230] <= 18'h21c50;
	 filter_out_expected[2231] <= 18'h14f48;
	 filter_out_expected[2232] <= 18'h37366;
	 filter_out_expected[2233] <= 18'h1c478;
	 filter_out_expected[2234] <= 18'h19e38;
	 filter_out_expected[2235] <= 18'h2f7e0;
	 filter_out_expected[2236] <= 18'h0c3b2;
	 filter_out_expected[2237] <= 18'h20afb;
	 filter_out_expected[2238] <= 18'h215b9;
	 filter_out_expected[2239] <= 18'h0b3c5;
	 filter_out_expected[2240] <= 18'h2ea85;
	 filter_out_expected[2241] <= 18'h2350c;
	 filter_out_expected[2242] <= 18'h31cbd;
	 filter_out_expected[2243] <= 18'h0a7cb;
	 filter_out_expected[2244] <= 18'h18d12;
	 filter_out_expected[2245] <= 18'h15757;
	 filter_out_expected[2246] <= 18'h0391f;
	 filter_out_expected[2247] <= 18'h324aa;
	 filter_out_expected[2248] <= 18'h2e868;
	 filter_out_expected[2249] <= 18'h35a41;
	 filter_out_expected[2250] <= 18'h3d4c4;
	 filter_out_expected[2251] <= 18'h039d7;
	 filter_out_expected[2252] <= 18'h08c6d;
	 filter_out_expected[2253] <= 18'h0865f;
	 filter_out_expected[2254] <= 18'h008d3;
	 filter_out_expected[2255] <= 18'h3bd27;
	 filter_out_expected[2256] <= 18'h3f781;
	 filter_out_expected[2257] <= 18'h0593a;
	 filter_out_expected[2258] <= 18'h07987;
	 filter_out_expected[2259] <= 18'h03023;
	 filter_out_expected[2260] <= 18'h3b997;
	 filter_out_expected[2261] <= 18'h35ebd;
	 filter_out_expected[2262] <= 18'h3536b;
	 filter_out_expected[2263] <= 18'h38a6c;
	 filter_out_expected[2264] <= 18'h3c641;
	 filter_out_expected[2265] <= 18'h3f65c;
	 filter_out_expected[2266] <= 18'h01ead;
	 filter_out_expected[2267] <= 18'h0572d;
	 filter_out_expected[2268] <= 18'h0d5cc;
	 filter_out_expected[2269] <= 18'h129b4;
	 filter_out_expected[2270] <= 18'h0f705;
	 filter_out_expected[2271] <= 18'h0607c;
	 filter_out_expected[2272] <= 18'h38ec1;
	 filter_out_expected[2273] <= 18'h2cb14;
	 filter_out_expected[2274] <= 18'h2a373;
	 filter_out_expected[2275] <= 18'h31099;
	 filter_out_expected[2276] <= 18'h3cf66;
	 filter_out_expected[2277] <= 18'h0ba40;
	 filter_out_expected[2278] <= 18'h1653d;
	 filter_out_expected[2279] <= 18'h14c1a;
	 filter_out_expected[2280] <= 18'h030de;
	 filter_out_expected[2281] <= 18'h2c89f;
	 filter_out_expected[2282] <= 18'h23993;
	 filter_out_expected[2283] <= 18'h2d100;
	 filter_out_expected[2284] <= 18'h01787;
	 filter_out_expected[2285] <= 18'h11cac;
	 filter_out_expected[2286] <= 18'h13cfb;
	 filter_out_expected[2287] <= 18'h0b9fd;
	 filter_out_expected[2288] <= 18'h00c9e;
	 filter_out_expected[2289] <= 18'h38344;
	 filter_out_expected[2290] <= 18'h34929;
	 filter_out_expected[2291] <= 18'h368a2;
	 filter_out_expected[2292] <= 18'h392e6;
	 filter_out_expected[2293] <= 18'h3e717;
	 filter_out_expected[2294] <= 18'h0624b;
	 filter_out_expected[2295] <= 18'h095e7;
	 filter_out_expected[2296] <= 18'h07151;
	 filter_out_expected[2297] <= 18'h02610;
	 filter_out_expected[2298] <= 18'h3ff04;
	 filter_out_expected[2299] <= 18'h00046;
	 filter_out_expected[2300] <= 18'h3f8ae;
	 filter_out_expected[2301] <= 18'h3d3a6;
	 filter_out_expected[2302] <= 18'h3bc5e;
	 filter_out_expected[2303] <= 18'h3d1c3;
	 filter_out_expected[2304] <= 18'h3f0df;
	 filter_out_expected[2305] <= 18'h03407;
	 filter_out_expected[2306] <= 18'h09cf5;
	 filter_out_expected[2307] <= 18'h0d037;
	 filter_out_expected[2308] <= 18'h03990;
	 filter_out_expected[2309] <= 18'h346ee;
	 filter_out_expected[2310] <= 18'h2faae;
	 filter_out_expected[2311] <= 18'h39e9f;
	 filter_out_expected[2312] <= 18'h0c47e;
	 filter_out_expected[2313] <= 18'h1692d;
	 filter_out_expected[2314] <= 18'h0dadb;
	 filter_out_expected[2315] <= 18'h39489;
	 filter_out_expected[2316] <= 18'h2e55d;
	 filter_out_expected[2317] <= 18'h343e4;
	 filter_out_expected[2318] <= 18'h3a91f;
	 filter_out_expected[2319] <= 18'h392e4;
	 filter_out_expected[2320] <= 18'h35ebb;
	 filter_out_expected[2321] <= 18'h3539d;
	 filter_out_expected[2322] <= 18'h3e688;
	 filter_out_expected[2323] <= 18'h0e8ea;
	 filter_out_expected[2324] <= 18'h16488;
	 filter_out_expected[2325] <= 18'h0a2a2;
	 filter_out_expected[2326] <= 18'h3454e;
	 filter_out_expected[2327] <= 18'h27e45;
	 filter_out_expected[2328] <= 18'h2d6fa;
	 filter_out_expected[2329] <= 18'h01210;
	 filter_out_expected[2330] <= 18'h17e3a;
	 filter_out_expected[2331] <= 18'h235fc;
	 filter_out_expected[2332] <= 18'h1d4c7;
	 filter_out_expected[2333] <= 18'h0a2a9;
	 filter_out_expected[2334] <= 18'h2f438;
	 filter_out_expected[2335] <= 18'h1722a;
	 filter_out_expected[2336] <= 18'h12d32;
	 filter_out_expected[2337] <= 18'h2c090;
	 filter_out_expected[2338] <= 18'h10242;
	 filter_out_expected[2339] <= 18'h1fa0c;
	 filter_out_expected[2340] <= 18'h15ceb;
	 filter_out_expected[2341] <= 18'h03ef1;
	 filter_out_expected[2342] <= 18'h37f32;
	 filter_out_expected[2343] <= 18'h36073;
	 filter_out_expected[2344] <= 18'h38449;
	 filter_out_expected[2345] <= 18'h3b875;
	 filter_out_expected[2346] <= 18'h02c8c;
	 filter_out_expected[2347] <= 18'h0d65e;
	 filter_out_expected[2348] <= 18'h15fda;
	 filter_out_expected[2349] <= 18'h1046e;
	 filter_out_expected[2350] <= 18'h3d311;
	 filter_out_expected[2351] <= 18'h2e87e;
	 filter_out_expected[2352] <= 18'h2f2d1;
	 filter_out_expected[2353] <= 18'h3cab9;
	 filter_out_expected[2354] <= 18'h0b7b3;
	 filter_out_expected[2355] <= 18'h0fba6;
	 filter_out_expected[2356] <= 18'h0450e;
	 filter_out_expected[2357] <= 18'h30627;
	 filter_out_expected[2358] <= 18'h22e7d;
	 filter_out_expected[2359] <= 18'h2b5b8;
	 filter_out_expected[2360] <= 18'h08246;
	 filter_out_expected[2361] <= 18'h217ef;
	 filter_out_expected[2362] <= 18'h223b9;
	 filter_out_expected[2363] <= 18'h07d91;
	 filter_out_expected[2364] <= 18'h24764;
	 filter_out_expected[2365] <= 18'h143ab;
	 filter_out_expected[2366] <= 18'h24032;
	 filter_out_expected[2367] <= 18'h0251f;
	 filter_out_expected[2368] <= 18'h1507f;
	 filter_out_expected[2369] <= 18'h130e5;
	 filter_out_expected[2370] <= 18'h051a5;
	 filter_out_expected[2371] <= 18'h3be79;
	 filter_out_expected[2372] <= 18'h3ea71;
	 filter_out_expected[2373] <= 18'h08773;
	 filter_out_expected[2374] <= 18'h11dfd;
	 filter_out_expected[2375] <= 18'h1489a;
	 filter_out_expected[2376] <= 18'h0e387;
	 filter_out_expected[2377] <= 18'h3e627;
	 filter_out_expected[2378] <= 18'h2d4e7;
	 filter_out_expected[2379] <= 18'h263af;
	 filter_out_expected[2380] <= 18'h290b8;
	 filter_out_expected[2381] <= 18'h306ef;
	 filter_out_expected[2382] <= 18'h3bfb9;
	 filter_out_expected[2383] <= 18'h09dfa;
	 filter_out_expected[2384] <= 18'h121a0;
	 filter_out_expected[2385] <= 18'h0f6e1;
	 filter_out_expected[2386] <= 18'h0288e;
	 filter_out_expected[2387] <= 18'h38b36;
	 filter_out_expected[2388] <= 18'h3df24;
	 filter_out_expected[2389] <= 18'h0ed36;
	 filter_out_expected[2390] <= 18'h19325;
	 filter_out_expected[2391] <= 18'h0e44d;
	 filter_out_expected[2392] <= 18'h333d6;
	 filter_out_expected[2393] <= 18'h1c201;
	 filter_out_expected[2394] <= 18'h1bf31;
	 filter_out_expected[2395] <= 18'h30665;
	 filter_out_expected[2396] <= 18'h0ab02;
	 filter_out_expected[2397] <= 18'h18ed2;
	 filter_out_expected[2398] <= 18'h116b7;
	 filter_out_expected[2399] <= 18'h3bd7d;
	 filter_out_expected[2400] <= 18'h30086;
	 filter_out_expected[2401] <= 18'h3cae0;
	 filter_out_expected[2402] <= 18'h14b30;
	 filter_out_expected[2403] <= 18'h1f599;
	 filter_out_expected[2404] <= 18'h0e760;
	 filter_out_expected[2405] <= 18'h2e8a2;
	 filter_out_expected[2406] <= 18'h1a94d;
	 filter_out_expected[2407] <= 18'h248bc;
	 filter_out_expected[2408] <= 18'h04913;
	 filter_out_expected[2409] <= 18'h1d909;
	 filter_out_expected[2410] <= 18'h1be85;
	 filter_out_expected[2411] <= 18'h09147;
	 filter_out_expected[2412] <= 18'h36ab8;
	 filter_out_expected[2413] <= 18'h2e055;
	 filter_out_expected[2414] <= 18'h2d3c3;
	 filter_out_expected[2415] <= 18'h32b42;
	 filter_out_expected[2416] <= 18'h3e402;
	 filter_out_expected[2417] <= 18'h0a674;
	 filter_out_expected[2418] <= 18'h12fa5;
	 filter_out_expected[2419] <= 18'h145a4;
	 filter_out_expected[2420] <= 18'h0cd2a;
	 filter_out_expected[2421] <= 18'h3f5ff;
	 filter_out_expected[2422] <= 18'h357ab;
	 filter_out_expected[2423] <= 18'h2edf6;
	 filter_out_expected[2424] <= 18'h29558;
	 filter_out_expected[2425] <= 18'h2c85c;
	 filter_out_expected[2426] <= 18'h3c237;
	 filter_out_expected[2427] <= 18'h0db54;
	 filter_out_expected[2428] <= 18'h11598;
	 filter_out_expected[2429] <= 18'h084ec;
	 filter_out_expected[2430] <= 18'h3d6a1;
	 filter_out_expected[2431] <= 18'h3bb84;
	 filter_out_expected[2432] <= 18'h0520c;
	 filter_out_expected[2433] <= 18'h0dc09;
	 filter_out_expected[2434] <= 18'h074ff;
	 filter_out_expected[2435] <= 18'h33a82;
	 filter_out_expected[2436] <= 18'h2bde7;
	 filter_out_expected[2437] <= 18'h3a544;
	 filter_out_expected[2438] <= 18'h0ea88;
	 filter_out_expected[2439] <= 18'h155a8;
	 filter_out_expected[2440] <= 18'h0c3e1;
	 filter_out_expected[2441] <= 18'h3cdaa;
	 filter_out_expected[2442] <= 18'h327bb;
	 filter_out_expected[2443] <= 18'h34d52;
	 filter_out_expected[2444] <= 18'h3de6a;
	 filter_out_expected[2445] <= 18'h04343;
	 filter_out_expected[2446] <= 18'h0317f;
	 filter_out_expected[2447] <= 18'h3d89c;
	 filter_out_expected[2448] <= 18'h36f25;
	 filter_out_expected[2449] <= 18'h3566e;
	 filter_out_expected[2450] <= 18'h3cdb1;
	 filter_out_expected[2451] <= 18'h0587d;
	 filter_out_expected[2452] <= 18'h02dea;
	 filter_out_expected[2453] <= 18'h36bf1;
	 filter_out_expected[2454] <= 18'h32cd3;
	 filter_out_expected[2455] <= 18'h3cc6c;
	 filter_out_expected[2456] <= 18'h0e2dc;
	 filter_out_expected[2457] <= 18'h1ce3c;
	 filter_out_expected[2458] <= 18'h20395;
	 filter_out_expected[2459] <= 18'h168aa;
	 filter_out_expected[2460] <= 18'h03a25;
	 filter_out_expected[2461] <= 18'h2f97b;
	 filter_out_expected[2462] <= 18'h24fe8;
	 filter_out_expected[2463] <= 18'h27553;
	 filter_out_expected[2464] <= 18'h32f94;
	 filter_out_expected[2465] <= 18'h01779;
	 filter_out_expected[2466] <= 18'h06444;
	 filter_out_expected[2467] <= 18'h3cf54;
	 filter_out_expected[2468] <= 18'h2d9fc;
	 filter_out_expected[2469] <= 18'h26649;
	 filter_out_expected[2470] <= 18'h2f028;
	 filter_out_expected[2471] <= 18'h0348f;
	 filter_out_expected[2472] <= 18'h18aec;
	 filter_out_expected[2473] <= 18'h2470e;
	 filter_out_expected[2474] <= 18'h207f5;
	 filter_out_expected[2475] <= 18'h10c99;
	 filter_out_expected[2476] <= 18'h02af8;
	 filter_out_expected[2477] <= 18'h37bd2;
	 filter_out_expected[2478] <= 18'h30b9b;
	 filter_out_expected[2479] <= 18'h31c4b;
	 filter_out_expected[2480] <= 18'h36b3e;
	 filter_out_expected[2481] <= 18'h39311;
	 filter_out_expected[2482] <= 18'h38e8d;
	 filter_out_expected[2483] <= 18'h396bf;
	 filter_out_expected[2484] <= 18'h39bfb;
	 filter_out_expected[2485] <= 18'h39927;
	 filter_out_expected[2486] <= 18'h3e6bc;
	 filter_out_expected[2487] <= 18'h0d7ad;
	 filter_out_expected[2488] <= 18'h1a053;
	 filter_out_expected[2489] <= 18'h16a29;
	 filter_out_expected[2490] <= 18'h0584f;
	 filter_out_expected[2491] <= 18'h31c3e;
	 filter_out_expected[2492] <= 18'h2a7bb;
	 filter_out_expected[2493] <= 18'h3360c;
	 filter_out_expected[2494] <= 18'h03b95;
	 filter_out_expected[2495] <= 18'h0f6a5;
	 filter_out_expected[2496] <= 18'h1002d;
	 filter_out_expected[2497] <= 18'h0616b;
	 filter_out_expected[2498] <= 18'h36870;
	 filter_out_expected[2499] <= 18'h292d5;
	 filter_out_expected[2500] <= 18'h2913d;
	 filter_out_expected[2501] <= 18'h3ae76;
	 filter_out_expected[2502] <= 18'h11225;
	 filter_out_expected[2503] <= 18'h198b6;
	 filter_out_expected[2504] <= 18'h124c5;
	 filter_out_expected[2505] <= 18'h062a5;
	 filter_out_expected[2506] <= 18'h3ab50;
	 filter_out_expected[2507] <= 18'h32e92;
	 filter_out_expected[2508] <= 18'h2f4dd;
	 filter_out_expected[2509] <= 18'h2fc88;
	 filter_out_expected[2510] <= 18'h37542;
	 filter_out_expected[2511] <= 18'h04886;
	 filter_out_expected[2512] <= 18'h11789;
	 filter_out_expected[2513] <= 18'h134b1;
	 filter_out_expected[2514] <= 18'h05ad7;
	 filter_out_expected[2515] <= 18'h358d8;
	 filter_out_expected[2516] <= 18'h2fc9d;
	 filter_out_expected[2517] <= 18'h341f5;
	 filter_out_expected[2518] <= 18'h3c103;
	 filter_out_expected[2519] <= 18'h00b45;
	 filter_out_expected[2520] <= 18'h05153;
	 filter_out_expected[2521] <= 18'h0fc43;
	 filter_out_expected[2522] <= 18'h18c0d;
	 filter_out_expected[2523] <= 18'h13ad5;
	 filter_out_expected[2524] <= 18'h02bd7;
	 filter_out_expected[2525] <= 18'h35445;
	 filter_out_expected[2526] <= 18'h32947;
	 filter_out_expected[2527] <= 18'h36fc6;
	 filter_out_expected[2528] <= 18'h3848c;
	 filter_out_expected[2529] <= 18'h35fd1;
	 filter_out_expected[2530] <= 18'h37587;
	 filter_out_expected[2531] <= 18'h3df86;
	 filter_out_expected[2532] <= 18'h06233;
	 filter_out_expected[2533] <= 18'h078f1;
	 filter_out_expected[2534] <= 18'h058b4;
	 filter_out_expected[2535] <= 18'h0408c;
	 filter_out_expected[2536] <= 18'h0027d;
	 filter_out_expected[2537] <= 18'h3ab9d;
	 filter_out_expected[2538] <= 18'h3dd01;
	 filter_out_expected[2539] <= 18'h095cd;
	 filter_out_expected[2540] <= 18'h12644;
	 filter_out_expected[2541] <= 18'h0e2f1;
	 filter_out_expected[2542] <= 18'h378af;
	 filter_out_expected[2543] <= 18'h1e489;
	 filter_out_expected[2544] <= 18'h172bf;
	 filter_out_expected[2545] <= 18'h27a84;
	 filter_out_expected[2546] <= 18'h048aa;
	 filter_out_expected[2547] <= 18'h1946e;
	 filter_out_expected[2548] <= 18'h1dad1;
	 filter_out_expected[2549] <= 18'h15ae5;
	 filter_out_expected[2550] <= 18'h09fb1;
	 filter_out_expected[2551] <= 18'h02629;
	 filter_out_expected[2552] <= 18'h3f1f3;
	 filter_out_expected[2553] <= 18'h3b560;
	 filter_out_expected[2554] <= 18'h3221a;
	 filter_out_expected[2555] <= 18'h27a38;
	 filter_out_expected[2556] <= 18'h2222f;
	 filter_out_expected[2557] <= 18'h2c614;
	 filter_out_expected[2558] <= 18'h0697f;
	 filter_out_expected[2559] <= 18'h24d2f;
	 filter_out_expected[2560] <= 18'h32d6d;
	 filter_out_expected[2561] <= 18'h21eb1;
	 filter_out_expected[2562] <= 18'h3be71;
	 filter_out_expected[2563] <= 18'h1f17c;
	 filter_out_expected[2564] <= 18'h1f4fe;
	 filter_out_expected[2565] <= 18'h32f63;
	 filter_out_expected[2566] <= 18'h08773;
	 filter_out_expected[2567] <= 18'h0d7ee;
	 filter_out_expected[2568] <= 18'h0154a;
	 filter_out_expected[2569] <= 18'h35295;
	 filter_out_expected[2570] <= 18'h3416c;
	 filter_out_expected[2571] <= 18'h3a645;
	 filter_out_expected[2572] <= 18'h02053;
	 filter_out_expected[2573] <= 18'h071e7;
	 filter_out_expected[2574] <= 18'h08f92;
	 filter_out_expected[2575] <= 18'h08212;
	 filter_out_expected[2576] <= 18'h04b2e;
	 filter_out_expected[2577] <= 18'h034a4;
	 filter_out_expected[2578] <= 18'h04ace;
	 filter_out_expected[2579] <= 18'h06510;
	 filter_out_expected[2580] <= 18'h02bbc;
	 filter_out_expected[2581] <= 18'h37d9b;
	 filter_out_expected[2582] <= 18'h3240c;
	 filter_out_expected[2583] <= 18'h3b138;
	 filter_out_expected[2584] <= 18'h0937d;
	 filter_out_expected[2585] <= 18'h0f089;
	 filter_out_expected[2586] <= 18'h048e7;
	 filter_out_expected[2587] <= 18'h30d85;
	 filter_out_expected[2588] <= 18'h28954;
	 filter_out_expected[2589] <= 18'h357c4;
	 filter_out_expected[2590] <= 18'h0b6b6;
	 filter_out_expected[2591] <= 18'h17764;
	 filter_out_expected[2592] <= 18'h1453a;
	 filter_out_expected[2593] <= 18'h07479;
	 filter_out_expected[2594] <= 18'h37d80;
	 filter_out_expected[2595] <= 18'h2f2b3;
	 filter_out_expected[2596] <= 18'h30313;
	 filter_out_expected[2597] <= 18'h373e0;
	 filter_out_expected[2598] <= 18'h3f488;
	 filter_out_expected[2599] <= 18'h01972;
	 filter_out_expected[2600] <= 18'h3d738;
	 filter_out_expected[2601] <= 18'h3908b;
	 filter_out_expected[2602] <= 18'h3ba47;
	 filter_out_expected[2603] <= 18'h06713;
	 filter_out_expected[2604] <= 18'h123eb;
	 filter_out_expected[2605] <= 18'h166f9;
	 filter_out_expected[2606] <= 18'h1023f;
	 filter_out_expected[2607] <= 18'h03aeb;
	 filter_out_expected[2608] <= 18'h383c8;
	 filter_out_expected[2609] <= 18'h32046;
	 filter_out_expected[2610] <= 18'h3056b;
	 filter_out_expected[2611] <= 18'h34f0f;
	 filter_out_expected[2612] <= 18'h39ce5;
	 filter_out_expected[2613] <= 18'h3776c;
	 filter_out_expected[2614] <= 18'h2e5a7;
	 filter_out_expected[2615] <= 18'h2b661;
	 filter_out_expected[2616] <= 18'h3aae3;
	 filter_out_expected[2617] <= 18'h14d0f;
	 filter_out_expected[2618] <= 18'h25da1;
	 filter_out_expected[2619] <= 18'h20237;
	 filter_out_expected[2620] <= 18'h0c7c0;
	 filter_out_expected[2621] <= 18'h3bcda;
	 filter_out_expected[2622] <= 18'h38041;
	 filter_out_expected[2623] <= 18'h3cf73;
	 filter_out_expected[2624] <= 18'h3bad7;
	 filter_out_expected[2625] <= 18'h30459;
	 filter_out_expected[2626] <= 18'h26109;
	 filter_out_expected[2627] <= 18'h26037;
	 filter_out_expected[2628] <= 18'h358fb;
	 filter_out_expected[2629] <= 18'h0e896;
	 filter_out_expected[2630] <= 18'h1e878;
	 filter_out_expected[2631] <= 18'h1926f;
	 filter_out_expected[2632] <= 18'h040be;
	 filter_out_expected[2633] <= 18'h352e3;
	 filter_out_expected[2634] <= 18'h387d8;
	 filter_out_expected[2635] <= 18'h045c8;
	 filter_out_expected[2636] <= 18'h0c025;
	 filter_out_expected[2637] <= 18'h062a3;
	 filter_out_expected[2638] <= 18'h34935;
	 filter_out_expected[2639] <= 18'h2a763;
	 filter_out_expected[2640] <= 18'h33011;
	 filter_out_expected[2641] <= 18'h051bb;
	 filter_out_expected[2642] <= 18'h100f6;
	 filter_out_expected[2643] <= 18'h08c99;
	 filter_out_expected[2644] <= 18'h37d70;
	 filter_out_expected[2645] <= 18'h30db5;
	 filter_out_expected[2646] <= 18'h3c68f;
	 filter_out_expected[2647] <= 18'h0f67c;
	 filter_out_expected[2648] <= 18'h134fc;
	 filter_out_expected[2649] <= 18'h07427;
	 filter_out_expected[2650] <= 18'h3e053;
	 filter_out_expected[2651] <= 18'h3e3d0;
	 filter_out_expected[2652] <= 18'h024a0;
	 filter_out_expected[2653] <= 18'h02cf1;
	 filter_out_expected[2654] <= 18'h00c58;
	 filter_out_expected[2655] <= 18'h007cf;
	 filter_out_expected[2656] <= 18'h01579;
	 filter_out_expected[2657] <= 18'h3c587;
	 filter_out_expected[2658] <= 18'h34d62;
	 filter_out_expected[2659] <= 18'h33701;
	 filter_out_expected[2660] <= 18'h3a844;
	 filter_out_expected[2661] <= 18'h04d51;
	 filter_out_expected[2662] <= 18'h0853e;
	 filter_out_expected[2663] <= 18'h06ef8;
	 filter_out_expected[2664] <= 18'h3ff8a;
	 filter_out_expected[2665] <= 18'h31b6b;
	 filter_out_expected[2666] <= 18'h23f52;
	 filter_out_expected[2667] <= 18'h23217;
	 filter_out_expected[2668] <= 18'h37fbe;
	 filter_out_expected[2669] <= 18'h1a607;
	 filter_out_expected[2670] <= 18'h31e11;
	 filter_out_expected[2671] <= 18'h2e34a;
	 filter_out_expected[2672] <= 18'h15048;
	 filter_out_expected[2673] <= 18'h35192;
	 filter_out_expected[2674] <= 18'h1dbc9;
	 filter_out_expected[2675] <= 18'h172c8;
	 filter_out_expected[2676] <= 18'h2272c;
	 filter_out_expected[2677] <= 18'h3b282;
	 filter_out_expected[2678] <= 18'h12a13;
	 filter_out_expected[2679] <= 18'h18f35;
	 filter_out_expected[2680] <= 18'h09cac;
	 filter_out_expected[2681] <= 18'h34377;
	 filter_out_expected[2682] <= 18'h2ce52;
	 filter_out_expected[2683] <= 18'h372fe;
	 filter_out_expected[2684] <= 18'h09af0;
	 filter_out_expected[2685] <= 18'h179dc;
	 filter_out_expected[2686] <= 18'h18453;
	 filter_out_expected[2687] <= 18'h0eaf5;
	 filter_out_expected[2688] <= 18'h04817;
	 filter_out_expected[2689] <= 18'h3e3a5;
	 filter_out_expected[2690] <= 18'h372ae;
	 filter_out_expected[2691] <= 18'h2df90;
	 filter_out_expected[2692] <= 18'h273a7;
	 filter_out_expected[2693] <= 18'h29a5d;
	 filter_out_expected[2694] <= 18'h3abda;
	 filter_out_expected[2695] <= 18'h11d9b;
	 filter_out_expected[2696] <= 18'h1b9a5;
	 filter_out_expected[2697] <= 18'h0c9c3;
	 filter_out_expected[2698] <= 18'h2fd89;
	 filter_out_expected[2699] <= 18'h1ed2c;
	 filter_out_expected[2700] <= 18'h2c693;
	 filter_out_expected[2701] <= 18'h0cf35;
	 filter_out_expected[2702] <= 18'h1fc5e;
	 filter_out_expected[2703] <= 18'h12484;
	 filter_out_expected[2704] <= 18'h36ba9;
	 filter_out_expected[2705] <= 18'h2e3ee;
	 filter_out_expected[2706] <= 18'h3d854;
	 filter_out_expected[2707] <= 18'h0fd37;
	 filter_out_expected[2708] <= 18'h0e044;
	 filter_out_expected[2709] <= 18'h39354;
	 filter_out_expected[2710] <= 18'h29eae;
	 filter_out_expected[2711] <= 18'h32692;
	 filter_out_expected[2712] <= 18'h0808e;
	 filter_out_expected[2713] <= 18'h16800;
	 filter_out_expected[2714] <= 18'h183ed;
	 filter_out_expected[2715] <= 18'h0e1ec;
	 filter_out_expected[2716] <= 18'h3c735;
	 filter_out_expected[2717] <= 18'h2b8e2;
	 filter_out_expected[2718] <= 18'h2394e;
	 filter_out_expected[2719] <= 18'h2a69c;
	 filter_out_expected[2720] <= 18'h3fb6a;
	 filter_out_expected[2721] <= 18'h163dd;
	 filter_out_expected[2722] <= 18'h1a0d0;
	 filter_out_expected[2723] <= 18'h07ef0;
	 filter_out_expected[2724] <= 18'h33f6b;
	 filter_out_expected[2725] <= 18'h324a9;
	 filter_out_expected[2726] <= 18'h3fe51;
	 filter_out_expected[2727] <= 18'h0cfe5;
	 filter_out_expected[2728] <= 18'h0e10e;
	 filter_out_expected[2729] <= 18'h004ea;
	 filter_out_expected[2730] <= 18'h34737;
	 filter_out_expected[2731] <= 18'h34f46;
	 filter_out_expected[2732] <= 18'h3c074;
	 filter_out_expected[2733] <= 18'h3f6a2;
	 filter_out_expected[2734] <= 18'h3a4f0;
	 filter_out_expected[2735] <= 18'h358a4;
	 filter_out_expected[2736] <= 18'h385b7;
	 filter_out_expected[2737] <= 18'h00d3e;
	 filter_out_expected[2738] <= 18'h0a1a1;
	 filter_out_expected[2739] <= 18'h10153;
	 filter_out_expected[2740] <= 18'h0b6d3;
	 filter_out_expected[2741] <= 18'h3f75b;
	 filter_out_expected[2742] <= 18'h34b6a;
	 filter_out_expected[2743] <= 18'h2ecef;
	 filter_out_expected[2744] <= 18'h2daea;
	 filter_out_expected[2745] <= 18'h3288e;
	 filter_out_expected[2746] <= 18'h03890;
	 filter_out_expected[2747] <= 18'h17a3f;
	 filter_out_expected[2748] <= 18'h1fb1c;
	 filter_out_expected[2749] <= 18'h154dd;
	 filter_out_expected[2750] <= 18'h3d54a;
	 filter_out_expected[2751] <= 18'h29618;
	 filter_out_expected[2752] <= 18'h2c92f;
	 filter_out_expected[2753] <= 18'h04b25;
	 filter_out_expected[2754] <= 18'h1a1e4;
	 filter_out_expected[2755] <= 18'h17fd9;
	 filter_out_expected[2756] <= 18'h3bf42;
	 filter_out_expected[2757] <= 18'h1c9de;
	 filter_out_expected[2758] <= 18'h1384c;
	 filter_out_expected[2759] <= 18'h2b988;
	 filter_out_expected[2760] <= 18'h124f0;
	 filter_out_expected[2761] <= 18'h25de0;
	 filter_out_expected[2762] <= 18'h1b35e;
	 filter_out_expected[2763] <= 18'h3fee0;
	 filter_out_expected[2764] <= 18'h2f524;
	 filter_out_expected[2765] <= 18'h3738c;
	 filter_out_expected[2766] <= 18'h09974;
	 filter_out_expected[2767] <= 18'h1357a;
	 filter_out_expected[2768] <= 18'h0bbdf;
	 filter_out_expected[2769] <= 18'h38333;
	 filter_out_expected[2770] <= 18'h28ebd;
	 filter_out_expected[2771] <= 18'h2743b;
	 filter_out_expected[2772] <= 18'h2e935;
	 filter_out_expected[2773] <= 18'h388a3;
	 filter_out_expected[2774] <= 18'h034ab;
	 filter_out_expected[2775] <= 18'h0ff14;
	 filter_out_expected[2776] <= 18'h189d7;
	 filter_out_expected[2777] <= 18'h1649f;
	 filter_out_expected[2778] <= 18'h0ef40;
	 filter_out_expected[2779] <= 18'h07418;
	 filter_out_expected[2780] <= 18'h3e981;
	 filter_out_expected[2781] <= 18'h328b4;
	 filter_out_expected[2782] <= 18'h2365c;
	 filter_out_expected[2783] <= 18'h1e02e;
	 filter_out_expected[2784] <= 18'h2f4f4;
	 filter_out_expected[2785] <= 18'h0cdcc;
	 filter_out_expected[2786] <= 18'h1a87b;
	 filter_out_expected[2787] <= 18'h0c3b4;
	 filter_out_expected[2788] <= 18'h384d8;
	 filter_out_expected[2789] <= 18'h3a792;
	 filter_out_expected[2790] <= 18'h0d11a;
	 filter_out_expected[2791] <= 18'h1569d;
	 filter_out_expected[2792] <= 18'h03c27;
	 filter_out_expected[2793] <= 18'h2b27b;
	 filter_out_expected[2794] <= 18'h294d6;
	 filter_out_expected[2795] <= 18'h3fae3;
	 filter_out_expected[2796] <= 18'h13583;
	 filter_out_expected[2797] <= 18'h10412;
	 filter_out_expected[2798] <= 18'h005b1;
	 filter_out_expected[2799] <= 18'h3686f;
	 filter_out_expected[2800] <= 18'h384e7;
	 filter_out_expected[2801] <= 18'h39b9e;
	 filter_out_expected[2802] <= 18'h38bcc;
	 filter_out_expected[2803] <= 18'h3cace;
	 filter_out_expected[2804] <= 18'h09fb6;
	 filter_out_expected[2805] <= 18'h14ba2;
	 filter_out_expected[2806] <= 18'h0cffb;
	 filter_out_expected[2807] <= 18'h391d3;
	 filter_out_expected[2808] <= 18'h2ec71;
	 filter_out_expected[2809] <= 18'h37b3a;
	 filter_out_expected[2810] <= 18'h02740;
	 filter_out_expected[2811] <= 18'h3ed8a;
	 filter_out_expected[2812] <= 18'h35345;
	 filter_out_expected[2813] <= 18'h3a74a;
	 filter_out_expected[2814] <= 18'h0b8f5;
	 filter_out_expected[2815] <= 18'h13595;
	 filter_out_expected[2816] <= 18'h07781;
	 filter_out_expected[2817] <= 18'h314e7;
	 filter_out_expected[2818] <= 18'h282f4;
	 filter_out_expected[2819] <= 18'h34ffd;
	 filter_out_expected[2820] <= 18'h0725a;
	 filter_out_expected[2821] <= 18'h09b65;
	 filter_out_expected[2822] <= 18'h00755;
	 filter_out_expected[2823] <= 18'h3d362;
	 filter_out_expected[2824] <= 18'h01058;
	 filter_out_expected[2825] <= 18'h05bcc;
	 filter_out_expected[2826] <= 18'h09ae6;
	 filter_out_expected[2827] <= 18'h0bd17;
	 filter_out_expected[2828] <= 18'h0985b;
	 filter_out_expected[2829] <= 18'h057e3;
	 filter_out_expected[2830] <= 18'h3f996;
	 filter_out_expected[2831] <= 18'h3256b;
	 filter_out_expected[2832] <= 18'h27ce2;
	 filter_out_expected[2833] <= 18'h2c7e4;
	 filter_out_expected[2834] <= 18'h3ed25;
	 filter_out_expected[2835] <= 18'h0dec9;
	 filter_out_expected[2836] <= 18'h0dbad;
	 filter_out_expected[2837] <= 18'h0223e;
	 filter_out_expected[2838] <= 18'h37321;
	 filter_out_expected[2839] <= 18'h3a324;
	 filter_out_expected[2840] <= 18'h05c32;
	 filter_out_expected[2841] <= 18'h0c537;
	 filter_out_expected[2842] <= 18'h0b6c0;
	 filter_out_expected[2843] <= 18'h09804;
	 filter_out_expected[2844] <= 18'h03cd7;
	 filter_out_expected[2845] <= 18'h39ef7;
	 filter_out_expected[2846] <= 18'h334c0;
	 filter_out_expected[2847] <= 18'h327eb;
	 filter_out_expected[2848] <= 18'h3c1df;
	 filter_out_expected[2849] <= 18'h06761;
	 filter_out_expected[2850] <= 18'h03a82;
	 filter_out_expected[2851] <= 18'h3719c;
	 filter_out_expected[2852] <= 18'h33a05;
	 filter_out_expected[2853] <= 18'h0279a;
	 filter_out_expected[2854] <= 18'h12734;
	 filter_out_expected[2855] <= 18'h0f43f;
	 filter_out_expected[2856] <= 18'h3a328;
	 filter_out_expected[2857] <= 18'h25824;
	 filter_out_expected[2858] <= 18'h22a07;
	 filter_out_expected[2859] <= 18'h39e10;
	 filter_out_expected[2860] <= 18'h169f2;
	 filter_out_expected[2861] <= 18'h1fd8f;
	 filter_out_expected[2862] <= 18'h17299;
	 filter_out_expected[2863] <= 18'h0ad63;
	 filter_out_expected[2864] <= 18'h01722;
	 filter_out_expected[2865] <= 18'h39549;
	 filter_out_expected[2866] <= 18'h30dd3;
	 filter_out_expected[2867] <= 18'h28933;
	 filter_out_expected[2868] <= 18'h25feb;
	 filter_out_expected[2869] <= 18'h2ffad;
	 filter_out_expected[2870] <= 18'h034c4;
	 filter_out_expected[2871] <= 18'h14cc5;
	 filter_out_expected[2872] <= 18'h2114e;
	 filter_out_expected[2873] <= 18'h255ff;
	 filter_out_expected[2874] <= 18'h190db;
	 filter_out_expected[2875] <= 18'h3c6f8;
	 filter_out_expected[2876] <= 18'h1efc2;
	 filter_out_expected[2877] <= 18'h12cb8;
	 filter_out_expected[2878] <= 18'h2037b;
	 filter_out_expected[2879] <= 18'h3da4e;
	 filter_out_expected[2880] <= 18'h1541a;
	 filter_out_expected[2881] <= 18'h19d81;
	 filter_out_expected[2882] <= 18'h0fb21;
	 filter_out_expected[2883] <= 18'h041cf;
	 filter_out_expected[2884] <= 18'h3e2e3;
	 filter_out_expected[2885] <= 18'h3d5f4;
	 filter_out_expected[2886] <= 18'h3ee13;
	 filter_out_expected[2887] <= 18'h3c4ef;
	 filter_out_expected[2888] <= 18'h3885c;
	 filter_out_expected[2889] <= 18'h3a336;
	 filter_out_expected[2890] <= 18'h01254;
	 filter_out_expected[2891] <= 18'h0805d;
	 filter_out_expected[2892] <= 18'h0a087;
	 filter_out_expected[2893] <= 18'h3fddf;
	 filter_out_expected[2894] <= 18'h2dfc8;
	 filter_out_expected[2895] <= 18'h26afc;
	 filter_out_expected[2896] <= 18'h33336;
	 filter_out_expected[2897] <= 18'h07d40;
	 filter_out_expected[2898] <= 18'h1042b;
	 filter_out_expected[2899] <= 18'h08469;
	 filter_out_expected[2900] <= 18'h39f8b;
	 filter_out_expected[2901] <= 18'h35d65;
	 filter_out_expected[2902] <= 18'h3f31d;
	 filter_out_expected[2903] <= 18'h08e17;
	 filter_out_expected[2904] <= 18'h07fc1;
	 filter_out_expected[2905] <= 18'h00e12;
	 filter_out_expected[2906] <= 18'h3bef8;
	 filter_out_expected[2907] <= 18'h3dcda;
	 filter_out_expected[2908] <= 18'h05977;
	 filter_out_expected[2909] <= 18'h0d516;
	 filter_out_expected[2910] <= 18'h0bfb6;
	 filter_out_expected[2911] <= 18'h3f0ee;
	 filter_out_expected[2912] <= 18'h33aac;
	 filter_out_expected[2913] <= 18'h3269f;
	 filter_out_expected[2914] <= 18'h38948;
	 filter_out_expected[2915] <= 18'h0106e;
	 filter_out_expected[2916] <= 18'h05d0a;
	 filter_out_expected[2917] <= 18'h07076;
	 filter_out_expected[2918] <= 18'h0cc82;
	 filter_out_expected[2919] <= 18'h16302;
	 filter_out_expected[2920] <= 18'h16f2f;
	 filter_out_expected[2921] <= 18'h06e0e;
	 filter_out_expected[2922] <= 18'h3127e;
	 filter_out_expected[2923] <= 18'h23b64;
	 filter_out_expected[2924] <= 18'h1fbd2;
	 filter_out_expected[2925] <= 18'h275de;
	 filter_out_expected[2926] <= 18'h3d3c5;
	 filter_out_expected[2927] <= 18'h16f2c;
	 filter_out_expected[2928] <= 18'h203f8;
	 filter_out_expected[2929] <= 18'h135b0;
	 filter_out_expected[2930] <= 18'h3d5d1;
	 filter_out_expected[2931] <= 18'h2d7b6;
	 filter_out_expected[2932] <= 18'h2a78e;
	 filter_out_expected[2933] <= 18'h302aa;
	 filter_out_expected[2934] <= 18'h35224;
	 filter_out_expected[2935] <= 18'h39263;
	 filter_out_expected[2936] <= 18'h062f0;
	 filter_out_expected[2937] <= 18'h19dc6;
	 filter_out_expected[2938] <= 18'h2356b;
	 filter_out_expected[2939] <= 18'h16655;
	 filter_out_expected[2940] <= 18'h3ae63;
	 filter_out_expected[2941] <= 18'h23586;
	 filter_out_expected[2942] <= 18'h189d4;
	 filter_out_expected[2943] <= 18'h1d768;
	 filter_out_expected[2944] <= 18'h2fdbc;
	 filter_out_expected[2945] <= 18'h0a87e;
	 filter_out_expected[2946] <= 18'h23d5b;
	 filter_out_expected[2947] <= 18'h2d83f;
	 filter_out_expected[2948] <= 18'h1dc2d;
	 filter_out_expected[2949] <= 18'h3df09;
	 filter_out_expected[2950] <= 18'h25a2e;
	 filter_out_expected[2951] <= 18'h24efd;
	 filter_out_expected[2952] <= 18'h336c8;
	 filter_out_expected[2953] <= 18'h00d6a;
	 filter_out_expected[2954] <= 18'h0666d;
	 filter_out_expected[2955] <= 18'h05708;
	 filter_out_expected[2956] <= 18'h055a8;
	 filter_out_expected[2957] <= 18'h04845;
	 filter_out_expected[2958] <= 18'h0024b;
	 filter_out_expected[2959] <= 18'h3df5e;
	 filter_out_expected[2960] <= 18'h03235;
	 filter_out_expected[2961] <= 18'h08309;
	 filter_out_expected[2962] <= 18'h04d9e;
	 filter_out_expected[2963] <= 18'h3a419;
	 filter_out_expected[2964] <= 18'h2fbef;
	 filter_out_expected[2965] <= 18'h2aa90;
	 filter_out_expected[2966] <= 18'h31a15;
	 filter_out_expected[2967] <= 18'h084ed;
	 filter_out_expected[2968] <= 18'h21a72;
	 filter_out_expected[2969] <= 18'h2a4ce;
	 filter_out_expected[2970] <= 18'h1a61b;
	 filter_out_expected[2971] <= 18'h3afb1;
	 filter_out_expected[2972] <= 18'h1e57c;
	 filter_out_expected[2973] <= 18'h16c54;
	 filter_out_expected[2974] <= 18'h258a8;
	 filter_out_expected[2975] <= 18'h3e50a;
	 filter_out_expected[2976] <= 18'h122fd;
	 filter_out_expected[2977] <= 18'h15b27;
	 filter_out_expected[2978] <= 18'h0a604;
	 filter_out_expected[2979] <= 18'h3c67e;
	 filter_out_expected[2980] <= 18'h347fa;
	 filter_out_expected[2981] <= 18'h38de0;
	 filter_out_expected[2982] <= 18'h047ea;
	 filter_out_expected[2983] <= 18'h05339;
	 filter_out_expected[2984] <= 18'h3b9ce;
	 filter_out_expected[2985] <= 18'h3a210;
	 filter_out_expected[2986] <= 18'h04be0;
	 filter_out_expected[2987] <= 18'h0acf0;
	 filter_out_expected[2988] <= 18'h019b8;
	 filter_out_expected[2989] <= 18'h32975;
	 filter_out_expected[2990] <= 18'h2f5a7;
	 filter_out_expected[2991] <= 18'h3bde7;
	 filter_out_expected[2992] <= 18'h10076;
	 filter_out_expected[2993] <= 18'h1aafa;
	 filter_out_expected[2994] <= 18'h12846;
	 filter_out_expected[2995] <= 18'h022a3;
	 filter_out_expected[2996] <= 18'h343ba;
	 filter_out_expected[2997] <= 18'h2bb91;
	 filter_out_expected[2998] <= 18'h28a22;
	 filter_out_expected[2999] <= 18'h328b1;
	 filter_out_expected[3000] <= 18'h04f2d;
	 filter_out_expected[3001] <= 18'h1239c;
	 filter_out_expected[3002] <= 18'h101f7;
	 filter_out_expected[3003] <= 18'h00e2b;
	 filter_out_expected[3004] <= 18'h33cbd;
	 filter_out_expected[3005] <= 18'h36017;
	 filter_out_expected[3006] <= 18'h06757;
	 filter_out_expected[3007] <= 18'h1386b;
	 filter_out_expected[3008] <= 18'h0ebc9;
	 filter_out_expected[3009] <= 18'h38fae;
	 filter_out_expected[3010] <= 18'h25f4e;
	 filter_out_expected[3011] <= 18'h258bb;
	 filter_out_expected[3012] <= 18'h397f4;
	 filter_out_expected[3013] <= 18'h11c50;
	 filter_out_expected[3014] <= 18'h1ce91;
	 filter_out_expected[3015] <= 18'h16257;
	 filter_out_expected[3016] <= 18'h0670f;
	 filter_out_expected[3017] <= 18'h3d60d;
	 filter_out_expected[3018] <= 18'h3c14d;
	 filter_out_expected[3019] <= 18'h3d4be;
	 filter_out_expected[3020] <= 18'h3ec65;
	 filter_out_expected[3021] <= 18'h3e69e;
	 filter_out_expected[3022] <= 18'h3b4aa;
	 filter_out_expected[3023] <= 18'h38846;
	 filter_out_expected[3024] <= 18'h37f7a;
	 filter_out_expected[3025] <= 18'h3adef;
	 filter_out_expected[3026] <= 18'h3df0d;
	 filter_out_expected[3027] <= 18'h3da1e;
	 filter_out_expected[3028] <= 18'h3e9df;
	 filter_out_expected[3029] <= 18'h02724;
	 filter_out_expected[3030] <= 18'h09762;
	 filter_out_expected[3031] <= 18'h0f5b8;
	 filter_out_expected[3032] <= 18'h073ca;
	 filter_out_expected[3033] <= 18'h35212;
	 filter_out_expected[3034] <= 18'h282dd;
	 filter_out_expected[3035] <= 18'h28274;
	 filter_out_expected[3036] <= 18'h32bc4;
	 filter_out_expected[3037] <= 18'h3e4fa;
	 filter_out_expected[3038] <= 18'h06fe3;
	 filter_out_expected[3039] <= 18'h10791;
	 filter_out_expected[3040] <= 18'h19c0f;
	 filter_out_expected[3041] <= 18'h1a8f3;
	 filter_out_expected[3042] <= 18'h0c4e3;
	 filter_out_expected[3043] <= 18'h32b2a;
	 filter_out_expected[3044] <= 18'h21882;
	 filter_out_expected[3045] <= 18'h28a7c;
	 filter_out_expected[3046] <= 18'h0020c;
	 filter_out_expected[3047] <= 18'h147df;
	 filter_out_expected[3048] <= 18'h180a1;
	 filter_out_expected[3049] <= 18'h0ca85;
	 filter_out_expected[3050] <= 18'h3d4d2;
	 filter_out_expected[3051] <= 18'h2fc1b;
	 filter_out_expected[3052] <= 18'h289b5;
	 filter_out_expected[3053] <= 18'h28645;
	 filter_out_expected[3054] <= 18'h32943;
	 filter_out_expected[3055] <= 18'h08b16;
	 filter_out_expected[3056] <= 18'h208d4;
	 filter_out_expected[3057] <= 18'h26e02;
	 filter_out_expected[3058] <= 18'h1319b;
	 filter_out_expected[3059] <= 18'h3308d;
	 filter_out_expected[3060] <= 18'h1ac0a;
	 filter_out_expected[3061] <= 18'h1919c;
	 filter_out_expected[3062] <= 18'h2d7a9;
	 filter_out_expected[3063] <= 18'h0f400;
	 filter_out_expected[3064] <= 18'h29ec6;
	 filter_out_expected[3065] <= 18'h2cebd;
	 filter_out_expected[3066] <= 18'h1926c;
	 filter_out_expected[3067] <= 18'h3ce2d;
	 filter_out_expected[3068] <= 18'h2a7bc;
	 filter_out_expected[3069] <= 18'h26d34;
	 filter_out_expected[3070] <= 18'h2a07d;
	 filter_out_expected[3071] <= 18'h2b6c8;
	 filter_out_expected[3072] <= 18'h2f8bf;
	 filter_out_expected[3073] <= 18'h3b9b7;
	 filter_out_expected[3074] <= 18'h0a610;
	 filter_out_expected[3075] <= 18'h0e7aa;
	 filter_out_expected[3076] <= 18'h03b58;
	 filter_out_expected[3077] <= 18'h39e37;
	 filter_out_expected[3078] <= 18'h3e733;
	 filter_out_expected[3079] <= 18'h0f610;
	 filter_out_expected[3080] <= 18'h19d1f;
	 filter_out_expected[3081] <= 18'h0f337;
	 filter_out_expected[3082] <= 18'h37b2b;
	 filter_out_expected[3083] <= 18'h2a5db;
	 filter_out_expected[3084] <= 18'h31049;
	 filter_out_expected[3085] <= 18'h0407b;
	 filter_out_expected[3086] <= 18'h13c09;
	 filter_out_expected[3087] <= 18'h104e3;
	 filter_out_expected[3088] <= 18'h3cb51;
	 filter_out_expected[3089] <= 18'h2a6ec;
	 filter_out_expected[3090] <= 18'h28c01;
	 filter_out_expected[3091] <= 18'h34092;
	 filter_out_expected[3092] <= 18'h026bb;
	 filter_out_expected[3093] <= 18'h0fed0;
	 filter_out_expected[3094] <= 18'h1a0eb;
	 filter_out_expected[3095] <= 18'h19497;
	 filter_out_expected[3096] <= 18'h0ca97;
	 filter_out_expected[3097] <= 18'h37b80;
	 filter_out_expected[3098] <= 18'h24364;
	 filter_out_expected[3099] <= 18'h22239;
	 filter_out_expected[3100] <= 18'h348f4;
	 filter_out_expected[3101] <= 18'h08dd1;
	 filter_out_expected[3102] <= 18'h0cf7d;
	 filter_out_expected[3103] <= 18'h05ff7;
	 filter_out_expected[3104] <= 18'h3b6c0;
	 filter_out_expected[3105] <= 18'h35019;
	 filter_out_expected[3106] <= 18'h3ac1f;
	 filter_out_expected[3107] <= 18'h0b43d;
	 filter_out_expected[3108] <= 18'h16c94;
	 filter_out_expected[3109] <= 18'h137ba;
	 filter_out_expected[3110] <= 18'h043d5;
	 filter_out_expected[3111] <= 18'h2fa68;
	 filter_out_expected[3112] <= 18'h20d84;
	 filter_out_expected[3113] <= 18'h2066c;
	 filter_out_expected[3114] <= 18'h2f17c;
	 filter_out_expected[3115] <= 18'h00ef6;
	 filter_out_expected[3116] <= 18'h11e20;
	 filter_out_expected[3117] <= 18'h1fd62;
	 filter_out_expected[3118] <= 18'h1d63a;
	 filter_out_expected[3119] <= 18'h0b3c5;
	 filter_out_expected[3120] <= 18'h366da;
	 filter_out_expected[3121] <= 18'h2b21f;
	 filter_out_expected[3122] <= 18'h2ab0e;
	 filter_out_expected[3123] <= 18'h337c2;
	 filter_out_expected[3124] <= 18'h00ac3;
	 filter_out_expected[3125] <= 18'h0c6ce;
	 filter_out_expected[3126] <= 18'h15378;
	 filter_out_expected[3127] <= 18'h18eef;
	 filter_out_expected[3128] <= 18'h126f7;
	 filter_out_expected[3129] <= 18'h3d5bb;
	 filter_out_expected[3130] <= 18'h297a7;
	 filter_out_expected[3131] <= 18'h25f15;
	 filter_out_expected[3132] <= 18'h30b22;
	 filter_out_expected[3133] <= 18'h3e86c;
	 filter_out_expected[3134] <= 18'h02a2b;
	 filter_out_expected[3135] <= 18'h3ef1c;
	 filter_out_expected[3136] <= 18'h3e76e;
	 filter_out_expected[3137] <= 18'h04e95;
	 filter_out_expected[3138] <= 18'h0bf5f;
	 filter_out_expected[3139] <= 18'h0bd79;
	 filter_out_expected[3140] <= 18'h058bf;
	 filter_out_expected[3141] <= 18'h00c6e;
	 filter_out_expected[3142] <= 18'h00f58;
	 filter_out_expected[3143] <= 18'h000ff;
	 filter_out_expected[3144] <= 18'h3c8ef;
	 filter_out_expected[3145] <= 18'h39ba9;
	 filter_out_expected[3146] <= 18'h3b391;
	 filter_out_expected[3147] <= 18'h3ef1e;
	 filter_out_expected[3148] <= 18'h00000;

	end // Input & Output data

endmodule
